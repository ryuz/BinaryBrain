`timescale 1ns / 1ps



module MnistStochasticLut6Mlp
        #(
            parameter USER_WIDTH = 0,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire                  reset,
            input  wire                  clk,
            input  wire                  cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [      784-1:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [       10-1:0]  out_data,
            output wire                  out_valid
        );


reg   [USER_BITS-1:0]  layer0_user;
wire  [     1024-1:0]  layer0_data;
reg                    layer0_valid;

MnistStochasticLut6Mlp_sub0
        #(
            .DEVICE     (DEVICE)
        )
    i_MnistStochasticLut6Mlp_sub0
        (
            .reset      (reset),
            .clk        (clk),
            .cke        (cke),
            
            .in_data    (in_data),
            .out_data   (layer0_data)
         );

always @(posedge clk) begin
    if ( reset ) begin
        layer0_user  <= {USER_BITS{1'bx}};
        layer0_valid <= 1'b0;
    end
    else if ( cke ) begin
        layer0_user  <= in_user;
        layer0_valid <= in_valid;
    end
end


reg   [USER_BITS-1:0]  layer1_user;
wire  [      360-1:0]  layer1_data;
reg                    layer1_valid;

MnistStochasticLut6Mlp_sub1
        #(
            .DEVICE     (DEVICE)
        )
    i_MnistStochasticLut6Mlp_sub1
        (
            .reset      (reset),
            .clk        (clk),
            .cke        (cke),
            
            .in_data    (layer0_data),
            .out_data   (layer1_data)
         );

always @(posedge clk) begin
    if ( reset ) begin
        layer1_user  <= {USER_BITS{1'bx}};
        layer1_valid <= 1'b0;
    end
    else if ( cke ) begin
        layer1_user  <= layer0_user;
        layer1_valid <= layer0_valid;
    end
end


reg   [USER_BITS-1:0]  layer2_user;
wire  [       60-1:0]  layer2_data;
reg                    layer2_valid;

MnistStochasticLut6Mlp_sub2
        #(
            .DEVICE     (DEVICE)
        )
    i_MnistStochasticLut6Mlp_sub2
        (
            .reset      (reset),
            .clk        (clk),
            .cke        (cke),
            
            .in_data    (layer1_data),
            .out_data   (layer2_data)
         );

always @(posedge clk) begin
    if ( reset ) begin
        layer2_user  <= {USER_BITS{1'bx}};
        layer2_valid <= 1'b0;
    end
    else if ( cke ) begin
        layer2_user  <= layer1_user;
        layer2_valid <= layer1_valid;
    end
end


reg   [USER_BITS-1:0]  layer3_user;
wire  [       10-1:0]  layer3_data;
reg                    layer3_valid;

MnistStochasticLut6Mlp_sub3
        #(
            .DEVICE     (DEVICE)
        )
    i_MnistStochasticLut6Mlp_sub3
        (
            .reset      (reset),
            .clk        (clk),
            .cke        (cke),
            
            .in_data    (layer2_data),
            .out_data   (layer3_data)
         );

always @(posedge clk) begin
    if ( reset ) begin
        layer3_user  <= {USER_BITS{1'bx}};
        layer3_valid <= 1'b0;
    end
    else if ( cke ) begin
        layer3_user  <= layer2_user;
        layer3_valid <= layer2_valid;
    end
end


assign out_data  = layer3_data;
assign out_user  = layer3_user;
assign out_valid = layer3_valid;

endmodule




module MnistStochasticLut6Mlp_sub0
        #(
            parameter DEVICE = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [783:0]  in_data,
            output wire [1023:0]  out_data
        );


// LUT : 0

wire lut_0_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111001101100001111110100001111001010101010100101010001010101),
            .DEVICE(DEVICE)
        )
    i_lut_0
        (
            .in_data({
                         in_data[111],
                         in_data[736],
                         in_data[420],
                         in_data[316],
                         in_data[302],
                         in_data[531]
                    }),
            .out_data(lut_0_out)
        );

reg   lut_0_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_0_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_0_ff <= lut_0_out;
    end
end

assign out_data[0] = lut_0_ff;




// LUT : 1

wire lut_1_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100100010010100110000111100110111101111101110000110001001100),
            .DEVICE(DEVICE)
        )
    i_lut_1
        (
            .in_data({
                         in_data[20],
                         in_data[400],
                         in_data[203],
                         in_data[529],
                         in_data[191],
                         in_data[73]
                    }),
            .out_data(lut_1_out)
        );

reg   lut_1_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1_ff <= lut_1_out;
    end
end

assign out_data[1] = lut_1_ff;




// LUT : 2

wire lut_2_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000110101111010011100111010110111010111011000111110101111110),
            .DEVICE(DEVICE)
        )
    i_lut_2
        (
            .in_data({
                         in_data[310],
                         in_data[148],
                         in_data[725],
                         in_data[692],
                         in_data[677],
                         in_data[620]
                    }),
            .out_data(lut_2_out)
        );

reg   lut_2_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_2_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_2_ff <= lut_2_out;
    end
end

assign out_data[2] = lut_2_ff;




// LUT : 3

wire lut_3_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000110011101010001001110000001011001011101111100110110111101100),
            .DEVICE(DEVICE)
        )
    i_lut_3
        (
            .in_data({
                         in_data[330],
                         in_data[606],
                         in_data[98],
                         in_data[501],
                         in_data[44],
                         in_data[663]
                    }),
            .out_data(lut_3_out)
        );

reg   lut_3_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_3_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_3_ff <= lut_3_out;
    end
end

assign out_data[3] = lut_3_ff;




// LUT : 4

wire lut_4_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001111111111000001110110010001101110010100000100111001000001010),
            .DEVICE(DEVICE)
        )
    i_lut_4
        (
            .in_data({
                         in_data[132],
                         in_data[707],
                         in_data[428],
                         in_data[129],
                         in_data[742],
                         in_data[334]
                    }),
            .out_data(lut_4_out)
        );

reg   lut_4_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_4_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_4_ff <= lut_4_out;
    end
end

assign out_data[4] = lut_4_ff;




// LUT : 5

wire lut_5_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110011101111101101111001010110110110000000000110111000011011),
            .DEVICE(DEVICE)
        )
    i_lut_5
        (
            .in_data({
                         in_data[574],
                         in_data[419],
                         in_data[699],
                         in_data[193],
                         in_data[298],
                         in_data[771]
                    }),
            .out_data(lut_5_out)
        );

reg   lut_5_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_5_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_5_ff <= lut_5_out;
    end
end

assign out_data[5] = lut_5_ff;




// LUT : 6

wire lut_6_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100001001000010001101110110001111000101000111100000110000001),
            .DEVICE(DEVICE)
        )
    i_lut_6
        (
            .in_data({
                         in_data[414],
                         in_data[359],
                         in_data[580],
                         in_data[40],
                         in_data[608],
                         in_data[783]
                    }),
            .out_data(lut_6_out)
        );

reg   lut_6_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_6_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_6_ff <= lut_6_out;
    end
end

assign out_data[6] = lut_6_ff;




// LUT : 7

wire lut_7_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100001111101011010101010100001100000001010011101100000000101),
            .DEVICE(DEVICE)
        )
    i_lut_7
        (
            .in_data({
                         in_data[338],
                         in_data[397],
                         in_data[424],
                         in_data[502],
                         in_data[320],
                         in_data[696]
                    }),
            .out_data(lut_7_out)
        );

reg   lut_7_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_7_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_7_ff <= lut_7_out;
    end
end

assign out_data[7] = lut_7_ff;




// LUT : 8

wire lut_8_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110110010010101001110011100000001000101000001010001010111000101),
            .DEVICE(DEVICE)
        )
    i_lut_8
        (
            .in_data({
                         in_data[394],
                         in_data[101],
                         in_data[512],
                         in_data[490],
                         in_data[480],
                         in_data[433]
                    }),
            .out_data(lut_8_out)
        );

reg   lut_8_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_8_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_8_ff <= lut_8_out;
    end
end

assign out_data[8] = lut_8_ff;




// LUT : 9

wire lut_9_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101000011101001001000100111100010011001110101111111110000110),
            .DEVICE(DEVICE)
        )
    i_lut_9
        (
            .in_data({
                         in_data[585],
                         in_data[322],
                         in_data[745],
                         in_data[472],
                         in_data[141],
                         in_data[355]
                    }),
            .out_data(lut_9_out)
        );

reg   lut_9_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_9_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_9_ff <= lut_9_out;
    end
end

assign out_data[9] = lut_9_ff;




// LUT : 10

wire lut_10_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010000100001011011001000000001100000010000110000111100110011),
            .DEVICE(DEVICE)
        )
    i_lut_10
        (
            .in_data({
                         in_data[561],
                         in_data[629],
                         in_data[252],
                         in_data[522],
                         in_data[753],
                         in_data[296]
                    }),
            .out_data(lut_10_out)
        );

reg   lut_10_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_10_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_10_ff <= lut_10_out;
    end
end

assign out_data[10] = lut_10_ff;




// LUT : 11

wire lut_11_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111111111101100001011101100110000100000100001001110000111101),
            .DEVICE(DEVICE)
        )
    i_lut_11
        (
            .in_data({
                         in_data[125],
                         in_data[426],
                         in_data[483],
                         in_data[560],
                         in_data[53],
                         in_data[689]
                    }),
            .out_data(lut_11_out)
        );

reg   lut_11_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_11_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_11_ff <= lut_11_out;
    end
end

assign out_data[11] = lut_11_ff;




// LUT : 12

wire lut_12_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011100001100000011111100100001111111000000000101101100000001),
            .DEVICE(DEVICE)
        )
    i_lut_12
        (
            .in_data({
                         in_data[123],
                         in_data[147],
                         in_data[340],
                         in_data[602],
                         in_data[171],
                         in_data[470]
                    }),
            .out_data(lut_12_out)
        );

reg   lut_12_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_12_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_12_ff <= lut_12_out;
    end
end

assign out_data[12] = lut_12_ff;




// LUT : 13

wire lut_13_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010100000000011111011110011101111110101110001110010010110000),
            .DEVICE(DEVICE)
        )
    i_lut_13
        (
            .in_data({
                         in_data[513],
                         in_data[690],
                         in_data[767],
                         in_data[168],
                         in_data[128],
                         in_data[232]
                    }),
            .out_data(lut_13_out)
        );

reg   lut_13_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_13_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_13_ff <= lut_13_out;
    end
end

assign out_data[13] = lut_13_ff;




// LUT : 14

wire lut_14_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001011111110101101011111001001101010111000111010011111101110001),
            .DEVICE(DEVICE)
        )
    i_lut_14
        (
            .in_data({
                         in_data[526],
                         in_data[276],
                         in_data[352],
                         in_data[104],
                         in_data[19],
                         in_data[94]
                    }),
            .out_data(lut_14_out)
        );

reg   lut_14_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_14_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_14_ff <= lut_14_out;
    end
end

assign out_data[14] = lut_14_ff;




// LUT : 15

wire lut_15_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001001110101100000101100101000000110001000000001100110000010),
            .DEVICE(DEVICE)
        )
    i_lut_15
        (
            .in_data({
                         in_data[600],
                         in_data[79],
                         in_data[267],
                         in_data[485],
                         in_data[446],
                         in_data[701]
                    }),
            .out_data(lut_15_out)
        );

reg   lut_15_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_15_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_15_ff <= lut_15_out;
    end
end

assign out_data[15] = lut_15_ff;




// LUT : 16

wire lut_16_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100110010010111110110101001010010000000010101000100111100111),
            .DEVICE(DEVICE)
        )
    i_lut_16
        (
            .in_data({
                         in_data[353],
                         in_data[116],
                         in_data[337],
                         in_data[58],
                         in_data[97],
                         in_data[368]
                    }),
            .out_data(lut_16_out)
        );

reg   lut_16_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_16_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_16_ff <= lut_16_out;
    end
end

assign out_data[16] = lut_16_ff;




// LUT : 17

wire lut_17_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001011110110100101111010011000100111100101011110110001011111111),
            .DEVICE(DEVICE)
        )
    i_lut_17
        (
            .in_data({
                         in_data[304],
                         in_data[221],
                         in_data[738],
                         in_data[481],
                         in_data[749],
                         in_data[77]
                    }),
            .out_data(lut_17_out)
        );

reg   lut_17_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_17_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_17_ff <= lut_17_out;
    end
end

assign out_data[17] = lut_17_ff;




// LUT : 18

wire lut_18_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111101010100110010001011010001100110100010100100101010101110),
            .DEVICE(DEVICE)
        )
    i_lut_18
        (
            .in_data({
                         in_data[152],
                         in_data[216],
                         in_data[33],
                         in_data[167],
                         in_data[374],
                         in_data[506]
                    }),
            .out_data(lut_18_out)
        );

reg   lut_18_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_18_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_18_ff <= lut_18_out;
    end
end

assign out_data[18] = lut_18_ff;




// LUT : 19

wire lut_19_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001101001011011001000110010001010000101001010100100010001000),
            .DEVICE(DEVICE)
        )
    i_lut_19
        (
            .in_data({
                         in_data[605],
                         in_data[389],
                         in_data[565],
                         in_data[728],
                         in_data[365],
                         in_data[166]
                    }),
            .out_data(lut_19_out)
        );

reg   lut_19_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_19_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_19_ff <= lut_19_out;
    end
end

assign out_data[19] = lut_19_ff;




// LUT : 20

wire lut_20_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011111011010001101010111000011110100110111000111000010111000),
            .DEVICE(DEVICE)
        )
    i_lut_20
        (
            .in_data({
                         in_data[64],
                         in_data[545],
                         in_data[436],
                         in_data[427],
                         in_data[172],
                         in_data[393]
                    }),
            .out_data(lut_20_out)
        );

reg   lut_20_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_20_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_20_ff <= lut_20_out;
    end
end

assign out_data[20] = lut_20_ff;




// LUT : 21

wire lut_21_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010011011010100001010000001100111100110101001111110011010100111),
            .DEVICE(DEVICE)
        )
    i_lut_21
        (
            .in_data({
                         in_data[54],
                         in_data[435],
                         in_data[549],
                         in_data[662],
                         in_data[26],
                         in_data[208]
                    }),
            .out_data(lut_21_out)
        );

reg   lut_21_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_21_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_21_ff <= lut_21_out;
    end
end

assign out_data[21] = lut_21_ff;




// LUT : 22

wire lut_22_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000011011110010000011100100111101010001011100000000000110011),
            .DEVICE(DEVICE)
        )
    i_lut_22
        (
            .in_data({
                         in_data[43],
                         in_data[107],
                         in_data[444],
                         in_data[628],
                         in_data[332],
                         in_data[431]
                    }),
            .out_data(lut_22_out)
        );

reg   lut_22_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_22_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_22_ff <= lut_22_out;
    end
end

assign out_data[22] = lut_22_ff;




// LUT : 23

wire lut_23_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000111101001000001100011101100101010000010000011001111110101),
            .DEVICE(DEVICE)
        )
    i_lut_23
        (
            .in_data({
                         in_data[648],
                         in_data[719],
                         in_data[195],
                         in_data[622],
                         in_data[489],
                         in_data[35]
                    }),
            .out_data(lut_23_out)
        );

reg   lut_23_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_23_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_23_ff <= lut_23_out;
    end
end

assign out_data[23] = lut_23_ff;




// LUT : 24

wire lut_24_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000000110000111100000111000010100101100000010001000010100000),
            .DEVICE(DEVICE)
        )
    i_lut_24
        (
            .in_data({
                         in_data[511],
                         in_data[155],
                         in_data[510],
                         in_data[724],
                         in_data[403],
                         in_data[269]
                    }),
            .out_data(lut_24_out)
        );

reg   lut_24_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_24_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_24_ff <= lut_24_out;
    end
end

assign out_data[24] = lut_24_ff;




// LUT : 25

wire lut_25_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010011011011000000010001001011100100101111101100101101111110),
            .DEVICE(DEVICE)
        )
    i_lut_25
        (
            .in_data({
                         in_data[63],
                         in_data[459],
                         in_data[504],
                         in_data[142],
                         in_data[176],
                         in_data[601]
                    }),
            .out_data(lut_25_out)
        );

reg   lut_25_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_25_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_25_ff <= lut_25_out;
    end
end

assign out_data[25] = lut_25_ff;




// LUT : 26

wire lut_26_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111111011101010101011111010010100000000000000010001100000010),
            .DEVICE(DEVICE)
        )
    i_lut_26
        (
            .in_data({
                         in_data[361],
                         in_data[236],
                         in_data[434],
                         in_data[718],
                         in_data[179],
                         in_data[131]
                    }),
            .out_data(lut_26_out)
        );

reg   lut_26_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_26_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_26_ff <= lut_26_out;
    end
end

assign out_data[26] = lut_26_ff;




// LUT : 27

wire lut_27_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000000001101000000001001000111000000001100000010000001000111),
            .DEVICE(DEVICE)
        )
    i_lut_27
        (
            .in_data({
                         in_data[717],
                         in_data[164],
                         in_data[494],
                         in_data[223],
                         in_data[521],
                         in_data[432]
                    }),
            .out_data(lut_27_out)
        );

reg   lut_27_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_27_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_27_ff <= lut_27_out;
    end
end

assign out_data[27] = lut_27_ff;




// LUT : 28

wire lut_28_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001011000111001100101101011010011100111011000101000110111101),
            .DEVICE(DEVICE)
        )
    i_lut_28
        (
            .in_data({
                         in_data[678],
                         in_data[774],
                         in_data[84],
                         in_data[634],
                         in_data[2],
                         in_data[528]
                    }),
            .out_data(lut_28_out)
        );

reg   lut_28_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_28_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_28_ff <= lut_28_out;
    end
end

assign out_data[28] = lut_28_ff;




// LUT : 29

wire lut_29_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001000011011110100010000100100101011100001101010001100001000),
            .DEVICE(DEVICE)
        )
    i_lut_29
        (
            .in_data({
                         in_data[706],
                         in_data[130],
                         in_data[186],
                         in_data[488],
                         in_data[42],
                         in_data[331]
                    }),
            .out_data(lut_29_out)
        );

reg   lut_29_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_29_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_29_ff <= lut_29_out;
    end
end

assign out_data[29] = lut_29_ff;




// LUT : 30

wire lut_30_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000001100000010000000100111101000001000010110011000100001110),
            .DEVICE(DEVICE)
        )
    i_lut_30
        (
            .in_data({
                         in_data[286],
                         in_data[99],
                         in_data[415],
                         in_data[333],
                         in_data[151],
                         in_data[576]
                    }),
            .out_data(lut_30_out)
        );

reg   lut_30_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_30_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_30_ff <= lut_30_out;
    end
end

assign out_data[30] = lut_30_ff;




// LUT : 31

wire lut_31_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101011100010101000101010010000110111011001111010010110000011),
            .DEVICE(DEVICE)
        )
    i_lut_31
        (
            .in_data({
                         in_data[228],
                         in_data[408],
                         in_data[160],
                         in_data[437],
                         in_data[779],
                         in_data[649]
                    }),
            .out_data(lut_31_out)
        );

reg   lut_31_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_31_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_31_ff <= lut_31_out;
    end
end

assign out_data[31] = lut_31_ff;




// LUT : 32

wire lut_32_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101011100100010110011110000001110000101100011011100000011000),
            .DEVICE(DEVICE)
        )
    i_lut_32
        (
            .in_data({
                         in_data[60],
                         in_data[465],
                         in_data[294],
                         in_data[402],
                         in_data[229],
                         in_data[587]
                    }),
            .out_data(lut_32_out)
        );

reg   lut_32_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_32_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_32_ff <= lut_32_out;
    end
end

assign out_data[32] = lut_32_ff;




// LUT : 33

wire lut_33_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001000101100011110011101110101110010011110101011000101010001),
            .DEVICE(DEVICE)
        )
    i_lut_33
        (
            .in_data({
                         in_data[396],
                         in_data[100],
                         in_data[318],
                         in_data[207],
                         in_data[204],
                         in_data[39]
                    }),
            .out_data(lut_33_out)
        );

reg   lut_33_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_33_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_33_ff <= lut_33_out;
    end
end

assign out_data[33] = lut_33_ff;




// LUT : 34

wire lut_34_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010111000101100100110000100011111010010101000100110011010011110),
            .DEVICE(DEVICE)
        )
    i_lut_34
        (
            .in_data({
                         in_data[292],
                         in_data[413],
                         in_data[76],
                         in_data[681],
                         in_data[756],
                         in_data[113]
                    }),
            .out_data(lut_34_out)
        );

reg   lut_34_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_34_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_34_ff <= lut_34_out;
    end
end

assign out_data[34] = lut_34_ff;




// LUT : 35

wire lut_35_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001101000110010100010010101001101100100001111101011101011110),
            .DEVICE(DEVICE)
        )
    i_lut_35
        (
            .in_data({
                         in_data[190],
                         in_data[14],
                         in_data[209],
                         in_data[418],
                         in_data[92],
                         in_data[590]
                    }),
            .out_data(lut_35_out)
        );

reg   lut_35_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_35_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_35_ff <= lut_35_out;
    end
end

assign out_data[35] = lut_35_ff;




// LUT : 36

wire lut_36_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001011000110101110100011110010111111111110111010101000111010000),
            .DEVICE(DEVICE)
        )
    i_lut_36
        (
            .in_data({
                         in_data[642],
                         in_data[652],
                         in_data[370],
                         in_data[367],
                         in_data[571],
                         in_data[727]
                    }),
            .out_data(lut_36_out)
        );

reg   lut_36_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_36_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_36_ff <= lut_36_out;
    end
end

assign out_data[36] = lut_36_ff;




// LUT : 37

wire lut_37_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100111001001011000000000100011110011010110011111011110110110),
            .DEVICE(DEVICE)
        )
    i_lut_37
        (
            .in_data({
                         in_data[22],
                         in_data[611],
                         in_data[482],
                         in_data[399],
                         in_data[478],
                         in_data[134]
                    }),
            .out_data(lut_37_out)
        );

reg   lut_37_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_37_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_37_ff <= lut_37_out;
    end
end

assign out_data[37] = lut_37_ff;




// LUT : 38

wire lut_38_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010000000000100100000000000000010000100010010001000000110001),
            .DEVICE(DEVICE)
        )
    i_lut_38
        (
            .in_data({
                         in_data[119],
                         in_data[429],
                         in_data[445],
                         in_data[491],
                         in_data[570],
                         in_data[487]
                    }),
            .out_data(lut_38_out)
        );

reg   lut_38_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_38_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_38_ff <= lut_38_out;
    end
end

assign out_data[38] = lut_38_ff;




// LUT : 39

wire lut_39_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110101110000110001100110110011001001101100000000000000010001110),
            .DEVICE(DEVICE)
        )
    i_lut_39
        (
            .in_data({
                         in_data[666],
                         in_data[215],
                         in_data[114],
                         in_data[404],
                         in_data[336],
                         in_data[328]
                    }),
            .out_data(lut_39_out)
        );

reg   lut_39_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_39_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_39_ff <= lut_39_out;
    end
end

assign out_data[39] = lut_39_ff;




// LUT : 40

wire lut_40_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100100101010000011000101011110101000011010100110111110110101),
            .DEVICE(DEVICE)
        )
    i_lut_40
        (
            .in_data({
                         in_data[364],
                         in_data[173],
                         in_data[326],
                         in_data[603],
                         in_data[5],
                         in_data[25]
                    }),
            .out_data(lut_40_out)
        );

reg   lut_40_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_40_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_40_ff <= lut_40_out;
    end
end

assign out_data[40] = lut_40_ff;




// LUT : 41

wire lut_41_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001011100110011111110101010001001001111111101111111101110000),
            .DEVICE(DEVICE)
        )
    i_lut_41
        (
            .in_data({
                         in_data[210],
                         in_data[452],
                         in_data[473],
                         in_data[462],
                         in_data[345],
                         in_data[174]
                    }),
            .out_data(lut_41_out)
        );

reg   lut_41_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_41_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_41_ff <= lut_41_out;
    end
end

assign out_data[41] = lut_41_ff;




// LUT : 42

wire lut_42_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001000101010101010101110101010010111101110100111111111111110),
            .DEVICE(DEVICE)
        )
    i_lut_42
        (
            .in_data({
                         in_data[238],
                         in_data[548],
                         in_data[598],
                         in_data[380],
                         in_data[635],
                         in_data[500]
                    }),
            .out_data(lut_42_out)
        );

reg   lut_42_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_42_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_42_ff <= lut_42_out;
    end
end

assign out_data[42] = lut_42_ff;




// LUT : 43

wire lut_43_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110010110100101111100010111000101010000110000000111101001111),
            .DEVICE(DEVICE)
        )
    i_lut_43
        (
            .in_data({
                         in_data[271],
                         in_data[138],
                         in_data[454],
                         in_data[307],
                         in_data[66],
                         in_data[91]
                    }),
            .out_data(lut_43_out)
        );

reg   lut_43_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_43_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_43_ff <= lut_43_out;
    end
end

assign out_data[43] = lut_43_ff;




// LUT : 44

wire lut_44_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001101001010100111101010111010011111101110011011101010001010100),
            .DEVICE(DEVICE)
        )
    i_lut_44
        (
            .in_data({
                         in_data[578],
                         in_data[672],
                         in_data[551],
                         in_data[640],
                         in_data[95],
                         in_data[137]
                    }),
            .out_data(lut_44_out)
        );

reg   lut_44_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_44_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_44_ff <= lut_44_out;
    end
end

assign out_data[44] = lut_44_ff;




// LUT : 45

wire lut_45_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001110000111101010101111100110010000101001011011101010100011100),
            .DEVICE(DEVICE)
        )
    i_lut_45
        (
            .in_data({
                         in_data[373],
                         in_data[451],
                         in_data[694],
                         in_data[671],
                         in_data[299],
                         in_data[460]
                    }),
            .out_data(lut_45_out)
        );

reg   lut_45_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_45_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_45_ff <= lut_45_out;
    end
end

assign out_data[45] = lut_45_ff;




// LUT : 46

wire lut_46_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001000011101000011011111010000000000001011001010111111111101),
            .DEVICE(DEVICE)
        )
    i_lut_46
        (
            .in_data({
                         in_data[509],
                         in_data[170],
                         in_data[750],
                         in_data[744],
                         in_data[261],
                         in_data[540]
                    }),
            .out_data(lut_46_out)
        );

reg   lut_46_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_46_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_46_ff <= lut_46_out;
    end
end

assign out_data[46] = lut_46_ff;




// LUT : 47

wire lut_47_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000011111100101010011111010101111011000000000010111011001110),
            .DEVICE(DEVICE)
        )
    i_lut_47
        (
            .in_data({
                         in_data[297],
                         in_data[70],
                         in_data[633],
                         in_data[288],
                         in_data[474],
                         in_data[83]
                    }),
            .out_data(lut_47_out)
        );

reg   lut_47_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_47_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_47_ff <= lut_47_out;
    end
end

assign out_data[47] = lut_47_ff;




// LUT : 48

wire lut_48_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111000010010101010101110011111010100010000101010100101110110),
            .DEVICE(DEVICE)
        )
    i_lut_48
        (
            .in_data({
                         in_data[751],
                         in_data[184],
                         in_data[117],
                         in_data[303],
                         in_data[245],
                         in_data[651]
                    }),
            .out_data(lut_48_out)
        );

reg   lut_48_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_48_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_48_ff <= lut_48_out;
    end
end

assign out_data[48] = lut_48_ff;




// LUT : 49

wire lut_49_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001010011100010110001011001011001110001111000100000001010100),
            .DEVICE(DEVICE)
        )
    i_lut_49
        (
            .in_data({
                         in_data[421],
                         in_data[375],
                         in_data[163],
                         in_data[664],
                         in_data[534],
                         in_data[56]
                    }),
            .out_data(lut_49_out)
        );

reg   lut_49_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_49_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_49_ff <= lut_49_out;
    end
end

assign out_data[49] = lut_49_ff;




// LUT : 50

wire lut_50_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110010101100000010000110000011000100000000010000000011110101),
            .DEVICE(DEVICE)
        )
    i_lut_50
        (
            .in_data({
                         in_data[306],
                         in_data[604],
                         in_data[277],
                         in_data[268],
                         in_data[458],
                         in_data[627]
                    }),
            .out_data(lut_50_out)
        );

reg   lut_50_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_50_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_50_ff <= lut_50_out;
    end
end

assign out_data[50] = lut_50_ff;




// LUT : 51

wire lut_51_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111011011001101100100001100110001101101010001000000000101010),
            .DEVICE(DEVICE)
        )
    i_lut_51
        (
            .in_data({
                         in_data[589],
                         in_data[213],
                         in_data[305],
                         in_data[547],
                         in_data[566],
                         in_data[740]
                    }),
            .out_data(lut_51_out)
        );

reg   lut_51_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_51_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_51_ff <= lut_51_out;
    end
end

assign out_data[51] = lut_51_ff;




// LUT : 52

wire lut_52_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011110000110010010001000001001111011001010011111110110100001),
            .DEVICE(DEVICE)
        )
    i_lut_52
        (
            .in_data({
                         in_data[165],
                         in_data[572],
                         in_data[126],
                         in_data[638],
                         in_data[31],
                         in_data[423]
                    }),
            .out_data(lut_52_out)
        );

reg   lut_52_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_52_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_52_ff <= lut_52_out;
    end
end

assign out_data[52] = lut_52_ff;




// LUT : 53

wire lut_53_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110100000010101110101101110101100101100011101010000011100010),
            .DEVICE(DEVICE)
        )
    i_lut_53
        (
            .in_data({
                         in_data[7],
                         in_data[667],
                         in_data[300],
                         in_data[564],
                         in_data[466],
                         in_data[192]
                    }),
            .out_data(lut_53_out)
        );

reg   lut_53_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_53_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_53_ff <= lut_53_out;
    end
end

assign out_data[53] = lut_53_ff;




// LUT : 54

wire lut_54_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101101001011010000000101000010111011001000011101100010001001),
            .DEVICE(DEVICE)
        )
    i_lut_54
        (
            .in_data({
                         in_data[23],
                         in_data[313],
                         in_data[543],
                         in_data[6],
                         in_data[537],
                         in_data[29]
                    }),
            .out_data(lut_54_out)
        );

reg   lut_54_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_54_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_54_ff <= lut_54_out;
    end
end

assign out_data[54] = lut_54_ff;




// LUT : 55

wire lut_55_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100110001001000000110000000000011111001101011100011011000011),
            .DEVICE(DEVICE)
        )
    i_lut_55
        (
            .in_data({
                         in_data[255],
                         in_data[15],
                         in_data[637],
                         in_data[527],
                         in_data[18],
                         in_data[467]
                    }),
            .out_data(lut_55_out)
        );

reg   lut_55_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_55_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_55_ff <= lut_55_out;
    end
end

assign out_data[55] = lut_55_ff;




// LUT : 56

wire lut_56_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000101111100111001000111000111111101000110010110100011000100),
            .DEVICE(DEVICE)
        )
    i_lut_56
        (
            .in_data({
                         in_data[729],
                         in_data[217],
                         in_data[106],
                         in_data[461],
                         in_data[759],
                         in_data[757]
                    }),
            .out_data(lut_56_out)
        );

reg   lut_56_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_56_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_56_ff <= lut_56_out;
    end
end

assign out_data[56] = lut_56_ff;




// LUT : 57

wire lut_57_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101001100011110110001100101011000000010001000100010001011011),
            .DEVICE(DEVICE)
        )
    i_lut_57
        (
            .in_data({
                         in_data[726],
                         in_data[146],
                         in_data[595],
                         in_data[242],
                         in_data[617],
                         in_data[650]
                    }),
            .out_data(lut_57_out)
        );

reg   lut_57_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_57_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_57_ff <= lut_57_out;
    end
end

assign out_data[57] = lut_57_ff;




// LUT : 58

wire lut_58_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010011011110010001001101000111111000101110001111000001111000),
            .DEVICE(DEVICE)
        )
    i_lut_58
        (
            .in_data({
                         in_data[395],
                         in_data[158],
                         in_data[350],
                         in_data[533],
                         in_data[463],
                         in_data[778]
                    }),
            .out_data(lut_58_out)
        );

reg   lut_58_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_58_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_58_ff <= lut_58_out;
    end
end

assign out_data[58] = lut_58_ff;




// LUT : 59

wire lut_59_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000110110101110110101010000000001011000000010001110010001110011),
            .DEVICE(DEVICE)
        )
    i_lut_59
        (
            .in_data({
                         in_data[655],
                         in_data[704],
                         in_data[746],
                         in_data[187],
                         in_data[777],
                         in_data[372]
                    }),
            .out_data(lut_59_out)
        );

reg   lut_59_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_59_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_59_ff <= lut_59_out;
    end
end

assign out_data[59] = lut_59_ff;




// LUT : 60

wire lut_60_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100111011101111010101000000110010011001111111011100101111111),
            .DEVICE(DEVICE)
        )
    i_lut_60
        (
            .in_data({
                         in_data[220],
                         in_data[703],
                         in_data[646],
                         in_data[665],
                         in_data[705],
                         in_data[291]
                    }),
            .out_data(lut_60_out)
        );

reg   lut_60_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_60_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_60_ff <= lut_60_out;
    end
end

assign out_data[60] = lut_60_ff;




// LUT : 61

wire lut_61_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001100100010101011010010111111101111000001001111101100001100),
            .DEVICE(DEVICE)
        )
    i_lut_61
        (
            .in_data({
                         in_data[630],
                         in_data[290],
                         in_data[96],
                         in_data[247],
                         in_data[136],
                         in_data[544]
                    }),
            .out_data(lut_61_out)
        );

reg   lut_61_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_61_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_61_ff <= lut_61_out;
    end
end

assign out_data[61] = lut_61_ff;




// LUT : 62

wire lut_62_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110001001101110001001101110111001100110011011100110111001101),
            .DEVICE(DEVICE)
        )
    i_lut_62
        (
            .in_data({
                         in_data[680],
                         in_data[497],
                         in_data[539],
                         in_data[360],
                         in_data[409],
                         in_data[455]
                    }),
            .out_data(lut_62_out)
        );

reg   lut_62_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_62_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_62_ff <= lut_62_out;
    end
end

assign out_data[62] = lut_62_ff;




// LUT : 63

wire lut_63_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011101010111010001000000010000010001100101110100111001011110010),
            .DEVICE(DEVICE)
        )
    i_lut_63
        (
            .in_data({
                         in_data[609],
                         in_data[686],
                         in_data[102],
                         in_data[175],
                         in_data[384],
                         in_data[591]
                    }),
            .out_data(lut_63_out)
        );

reg   lut_63_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_63_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_63_ff <= lut_63_out;
    end
end

assign out_data[63] = lut_63_ff;




// LUT : 64

wire lut_64_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100001101110100101010000010111110010110000100001101001110010011),
            .DEVICE(DEVICE)
        )
    i_lut_64
        (
            .in_data({
                         in_data[45],
                         in_data[448],
                         in_data[457],
                         in_data[89],
                         in_data[619],
                         in_data[382]
                    }),
            .out_data(lut_64_out)
        );

reg   lut_64_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_64_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_64_ff <= lut_64_out;
    end
end

assign out_data[64] = lut_64_ff;




// LUT : 65

wire lut_65_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001011100100011011100110111001100111100000001001111010001010),
            .DEVICE(DEVICE)
        )
    i_lut_65
        (
            .in_data({
                         in_data[185],
                         in_data[200],
                         in_data[21],
                         in_data[499],
                         in_data[162],
                         in_data[249]
                    }),
            .out_data(lut_65_out)
        );

reg   lut_65_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_65_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_65_ff <= lut_65_out;
    end
end

assign out_data[65] = lut_65_ff;




// LUT : 66

wire lut_66_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101010000011111010001010100010001000100000010110010111010101),
            .DEVICE(DEVICE)
        )
    i_lut_66
        (
            .in_data({
                         in_data[13],
                         in_data[573],
                         in_data[323],
                         in_data[122],
                         in_data[568],
                         in_data[765]
                    }),
            .out_data(lut_66_out)
        );

reg   lut_66_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_66_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_66_ff <= lut_66_out;
    end
end

assign out_data[66] = lut_66_ff;




// LUT : 67

wire lut_67_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000011001100000111101111111010001100100100011101111101001110),
            .DEVICE(DEVICE)
        )
    i_lut_67
        (
            .in_data({
                         in_data[214],
                         in_data[391],
                         in_data[410],
                         in_data[28],
                         in_data[149],
                         in_data[695]
                    }),
            .out_data(lut_67_out)
        );

reg   lut_67_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_67_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_67_ff <= lut_67_out;
    end
end

assign out_data[67] = lut_67_ff;




// LUT : 68

wire lut_68_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000110001100001100000010100111111100000010100110100001000100),
            .DEVICE(DEVICE)
        )
    i_lut_68
        (
            .in_data({
                         in_data[586],
                         in_data[782],
                         in_data[109],
                         in_data[516],
                         in_data[260],
                         in_data[67]
                    }),
            .out_data(lut_68_out)
        );

reg   lut_68_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_68_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_68_ff <= lut_68_out;
    end
end

assign out_data[68] = lut_68_ff;




// LUT : 69

wire lut_69_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111100000110001000110011011010101111000011100100111100100000),
            .DEVICE(DEVICE)
        )
    i_lut_69
        (
            .in_data({
                         in_data[65],
                         in_data[709],
                         in_data[441],
                         in_data[309],
                         in_data[284],
                         in_data[206]
                    }),
            .out_data(lut_69_out)
        );

reg   lut_69_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_69_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_69_ff <= lut_69_out;
    end
end

assign out_data[69] = lut_69_ff;




// LUT : 70

wire lut_70_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100011000010010000001101001011101010010000000111111011111111),
            .DEVICE(DEVICE)
        )
    i_lut_70
        (
            .in_data({
                         in_data[658],
                         in_data[582],
                         in_data[581],
                         in_data[327],
                         in_data[439],
                         in_data[280]
                    }),
            .out_data(lut_70_out)
        );

reg   lut_70_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_70_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_70_ff <= lut_70_out;
    end
end

assign out_data[70] = lut_70_ff;




// LUT : 71

wire lut_71_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100110111001110110100101011110100111000101110100001000001001),
            .DEVICE(DEVICE)
        )
    i_lut_71
        (
            .in_data({
                         in_data[623],
                         in_data[684],
                         in_data[530],
                         in_data[764],
                         in_data[732],
                         in_data[758]
                    }),
            .out_data(lut_71_out)
        );

reg   lut_71_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_71_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_71_ff <= lut_71_out;
    end
end

assign out_data[71] = lut_71_ff;




// LUT : 72

wire lut_72_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111101111101010111110111011111111111000100001111110100110010),
            .DEVICE(DEVICE)
        )
    i_lut_72
        (
            .in_data({
                         in_data[536],
                         in_data[262],
                         in_data[507],
                         in_data[324],
                         in_data[484],
                         in_data[86]
                    }),
            .out_data(lut_72_out)
        );

reg   lut_72_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_72_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_72_ff <= lut_72_out;
    end
end

assign out_data[72] = lut_72_ff;




// LUT : 73

wire lut_73_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100010101000110001111111000010100111010110001111001001011010),
            .DEVICE(DEVICE)
        )
    i_lut_73
        (
            .in_data({
                         in_data[82],
                         in_data[339],
                         in_data[234],
                         in_data[105],
                         in_data[246],
                         in_data[776]
                    }),
            .out_data(lut_73_out)
        );

reg   lut_73_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_73_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_73_ff <= lut_73_out;
    end
end

assign out_data[73] = lut_73_ff;




// LUT : 74

wire lut_74_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010011111110010111111100110010111111000110010011011101111111),
            .DEVICE(DEVICE)
        )
    i_lut_74
        (
            .in_data({
                         in_data[583],
                         in_data[254],
                         in_data[335],
                         in_data[317],
                         in_data[169],
                         in_data[702]
                    }),
            .out_data(lut_74_out)
        );

reg   lut_74_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_74_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_74_ff <= lut_74_out;
    end
end

assign out_data[74] = lut_74_ff;




// LUT : 75

wire lut_75_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001111100101001001101001010101000111111000101010101011010011),
            .DEVICE(DEVICE)
        )
    i_lut_75
        (
            .in_data({
                         in_data[201],
                         in_data[440],
                         in_data[256],
                         in_data[775],
                         in_data[59],
                         in_data[0]
                    }),
            .out_data(lut_75_out)
        );

reg   lut_75_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_75_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_75_ff <= lut_75_out;
    end
end

assign out_data[75] = lut_75_ff;




// LUT : 76

wire lut_76_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010111010101011010011101111100000100010111000000110001011111),
            .DEVICE(DEVICE)
        )
    i_lut_76
        (
            .in_data({
                         in_data[610],
                         in_data[401],
                         in_data[69],
                         in_data[358],
                         in_data[639],
                         in_data[406]
                    }),
            .out_data(lut_76_out)
        );

reg   lut_76_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_76_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_76_ff <= lut_76_out;
    end
end

assign out_data[76] = lut_76_ff;




// LUT : 77

wire lut_77_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001100110110000110101001111010101101110111101110010010101011000),
            .DEVICE(DEVICE)
        )
    i_lut_77
        (
            .in_data({
                         in_data[196],
                         in_data[281],
                         in_data[62],
                         in_data[673],
                         in_data[325],
                         in_data[739]
                    }),
            .out_data(lut_77_out)
        );

reg   lut_77_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_77_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_77_ff <= lut_77_out;
    end
end

assign out_data[77] = lut_77_ff;




// LUT : 78

wire lut_78_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111010011000000001100000001011001100110001100110110011100100),
            .DEVICE(DEVICE)
        )
    i_lut_78
        (
            .in_data({
                         in_data[225],
                         in_data[653],
                         in_data[579],
                         in_data[369],
                         in_data[405],
                         in_data[12]
                    }),
            .out_data(lut_78_out)
        );

reg   lut_78_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_78_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_78_ff <= lut_78_out;
    end
end

assign out_data[78] = lut_78_ff;




// LUT : 79

wire lut_79_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001111011111010100000001000010110001101101010001001100010011),
            .DEVICE(DEVICE)
        )
    i_lut_79
        (
            .in_data({
                         in_data[212],
                         in_data[593],
                         in_data[492],
                         in_data[257],
                         in_data[720],
                         in_data[180]
                    }),
            .out_data(lut_79_out)
        );

reg   lut_79_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_79_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_79_ff <= lut_79_out;
    end
end

assign out_data[79] = lut_79_ff;




// LUT : 80

wire lut_80_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111010001000000000001010001011000011111010101011110010110011),
            .DEVICE(DEVICE)
        )
    i_lut_80
        (
            .in_data({
                         in_data[520],
                         in_data[741],
                         in_data[670],
                         in_data[381],
                         in_data[773],
                         in_data[387]
                    }),
            .out_data(lut_80_out)
        );

reg   lut_80_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_80_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_80_ff <= lut_80_out;
    end
end

assign out_data[80] = lut_80_ff;




// LUT : 81

wire lut_81_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000001011100101010010111001101101100111010100000100111011110),
            .DEVICE(DEVICE)
        )
    i_lut_81
        (
            .in_data({
                         in_data[183],
                         in_data[710],
                         in_data[49],
                         in_data[390],
                         in_data[108],
                         in_data[584]
                    }),
            .out_data(lut_81_out)
        );

reg   lut_81_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_81_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_81_ff <= lut_81_out;
    end
end

assign out_data[81] = lut_81_ff;




// LUT : 82

wire lut_82_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110110111110011110111101000011100100110111110110000011100000000),
            .DEVICE(DEVICE)
        )
    i_lut_82
        (
            .in_data({
                         in_data[222],
                         in_data[514],
                         in_data[11],
                         in_data[453],
                         in_data[693],
                         in_data[265]
                    }),
            .out_data(lut_82_out)
        );

reg   lut_82_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_82_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_82_ff <= lut_82_out;
    end
end

assign out_data[82] = lut_82_ff;




// LUT : 83

wire lut_83_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101100011111001001001110101101010100001000001010111010001010),
            .DEVICE(DEVICE)
        )
    i_lut_83
        (
            .in_data({
                         in_data[647],
                         in_data[733],
                         in_data[178],
                         in_data[379],
                         in_data[293],
                         in_data[714]
                    }),
            .out_data(lut_83_out)
        );

reg   lut_83_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_83_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_83_ff <= lut_83_out;
    end
end

assign out_data[83] = lut_83_ff;




// LUT : 84

wire lut_84_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111011011111000111000001110000011111110111110011011111111100),
            .DEVICE(DEVICE)
        )
    i_lut_84
        (
            .in_data({
                         in_data[721],
                         in_data[592],
                         in_data[311],
                         in_data[442],
                         in_data[93],
                         in_data[518]
                    }),
            .out_data(lut_84_out)
        );

reg   lut_84_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_84_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_84_ff <= lut_84_out;
    end
end

assign out_data[84] = lut_84_ff;




// LUT : 85

wire lut_85_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010100010000010011111101001111111000001000010111000010111101),
            .DEVICE(DEVICE)
        )
    i_lut_85
        (
            .in_data({
                         in_data[4],
                         in_data[386],
                         in_data[181],
                         in_data[523],
                         in_data[17],
                         in_data[270]
                    }),
            .out_data(lut_85_out)
        );

reg   lut_85_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_85_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_85_ff <= lut_85_out;
    end
end

assign out_data[85] = lut_85_ff;




// LUT : 86

wire lut_86_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000101110101111100001111010001110100010101010111110111111111),
            .DEVICE(DEVICE)
        )
    i_lut_86
        (
            .in_data({
                         in_data[398],
                         in_data[272],
                         in_data[486],
                         in_data[535],
                         in_data[68],
                         in_data[351]
                    }),
            .out_data(lut_86_out)
        );

reg   lut_86_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_86_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_86_ff <= lut_86_out;
    end
end

assign out_data[86] = lut_86_ff;




// LUT : 87

wire lut_87_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001100110110010001100111011001101000101010010010011001000110),
            .DEVICE(DEVICE)
        )
    i_lut_87
        (
            .in_data({
                         in_data[713],
                         in_data[392],
                         in_data[577],
                         in_data[575],
                         in_data[371],
                         in_data[37]
                    }),
            .out_data(lut_87_out)
        );

reg   lut_87_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_87_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_87_ff <= lut_87_out;
    end
end

assign out_data[87] = lut_87_ff;




// LUT : 88

wire lut_88_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110011101100011100011001100111100010100010000000100111100001),
            .DEVICE(DEVICE)
        )
    i_lut_88
        (
            .in_data({
                         in_data[343],
                         in_data[243],
                         in_data[607],
                         in_data[538],
                         in_data[754],
                         in_data[283]
                    }),
            .out_data(lut_88_out)
        );

reg   lut_88_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_88_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_88_ff <= lut_88_out;
    end
end

assign out_data[88] = lut_88_ff;




// LUT : 89

wire lut_89_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110110000100001011001010110010101111000111111101000011100100),
            .DEVICE(DEVICE)
        )
    i_lut_89
        (
            .in_data({
                         in_data[161],
                         in_data[251],
                         in_data[626],
                         in_data[3],
                         in_data[687],
                         in_data[624]
                    }),
            .out_data(lut_89_out)
        );

reg   lut_89_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_89_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_89_ff <= lut_89_out;
    end
end

assign out_data[89] = lut_89_ff;




// LUT : 90

wire lut_90_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011010100010100000101010001000110110100101010001011100100010),
            .DEVICE(DEVICE)
        )
    i_lut_90
        (
            .in_data({
                         in_data[266],
                         in_data[237],
                         in_data[239],
                         in_data[295],
                         in_data[377],
                         in_data[674]
                    }),
            .out_data(lut_90_out)
        );

reg   lut_90_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_90_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_90_ff <= lut_90_out;
    end
end

assign out_data[90] = lut_90_ff;




// LUT : 91

wire lut_91_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001101100111001101101101111111011111011101101110011001011111110),
            .DEVICE(DEVICE)
        )
    i_lut_91
        (
            .in_data({
                         in_data[301],
                         in_data[231],
                         in_data[211],
                         in_data[596],
                         in_data[475],
                         in_data[417]
                    }),
            .out_data(lut_91_out)
        );

reg   lut_91_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_91_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_91_ff <= lut_91_out;
    end
end

assign out_data[91] = lut_91_ff;




// LUT : 92

wire lut_92_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100101000011011100011011010001001010010011111110111111111101),
            .DEVICE(DEVICE)
        )
    i_lut_92
        (
            .in_data({
                         in_data[1],
                         in_data[61],
                         in_data[139],
                         in_data[508],
                         in_data[41],
                         in_data[342]
                    }),
            .out_data(lut_92_out)
        );

reg   lut_92_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_92_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_92_ff <= lut_92_out;
    end
end

assign out_data[92] = lut_92_ff;




// LUT : 93

wire lut_93_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011110111100001100001001000000000101111111111001110010110001110),
            .DEVICE(DEVICE)
        )
    i_lut_93
        (
            .in_data({
                         in_data[55],
                         in_data[770],
                         in_data[218],
                         in_data[471],
                         in_data[226],
                         in_data[110]
                    }),
            .out_data(lut_93_out)
        );

reg   lut_93_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_93_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_93_ff <= lut_93_out;
    end
end

assign out_data[93] = lut_93_ff;




// LUT : 94

wire lut_94_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110110111001101011011110001011001111001100110011000100000000001),
            .DEVICE(DEVICE)
        )
    i_lut_94
        (
            .in_data({
                         in_data[422],
                         in_data[341],
                         in_data[781],
                         in_data[143],
                         in_data[616],
                         in_data[554]
                    }),
            .out_data(lut_94_out)
        );

reg   lut_94_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_94_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_94_ff <= lut_94_out;
    end
end

assign out_data[94] = lut_94_ff;




// LUT : 95

wire lut_95_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010011010010111110001100110000111000100011010111010001111011),
            .DEVICE(DEVICE)
        )
    i_lut_95
        (
            .in_data({
                         in_data[679],
                         in_data[731],
                         in_data[289],
                         in_data[154],
                         in_data[449],
                         in_data[456]
                    }),
            .out_data(lut_95_out)
        );

reg   lut_95_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_95_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_95_ff <= lut_95_out;
    end
end

assign out_data[95] = lut_95_ff;




// LUT : 96

wire lut_96_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111011111101000010101111111101011010110011000110001111111101),
            .DEVICE(DEVICE)
        )
    i_lut_96
        (
            .in_data({
                         in_data[552],
                         in_data[347],
                         in_data[32],
                         in_data[150],
                         in_data[632],
                         in_data[321]
                    }),
            .out_data(lut_96_out)
        );

reg   lut_96_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_96_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_96_ff <= lut_96_out;
    end
end

assign out_data[96] = lut_96_ff;




// LUT : 97

wire lut_97_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100001000101000101111001011101101101100110000000000000010111011),
            .DEVICE(DEVICE)
        )
    i_lut_97
        (
            .in_data({
                         in_data[416],
                         in_data[279],
                         in_data[378],
                         in_data[495],
                         in_data[762],
                         in_data[657]
                    }),
            .out_data(lut_97_out)
        );

reg   lut_97_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_97_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_97_ff <= lut_97_out;
    end
end

assign out_data[97] = lut_97_ff;




// LUT : 98

wire lut_98_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111110000011100011111110010111111010011010110011110011110101011),
            .DEVICE(DEVICE)
        )
    i_lut_98
        (
            .in_data({
                         in_data[362],
                         in_data[614],
                         in_data[524],
                         in_data[314],
                         in_data[219],
                         in_data[71]
                    }),
            .out_data(lut_98_out)
        );

reg   lut_98_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_98_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_98_ff <= lut_98_out;
    end
end

assign out_data[98] = lut_98_ff;




// LUT : 99

wire lut_99_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101100101011110110000011101100101100000101010000111110001010),
            .DEVICE(DEVICE)
        )
    i_lut_99
        (
            .in_data({
                         in_data[388],
                         in_data[763],
                         in_data[51],
                         in_data[755],
                         in_data[156],
                         in_data[75]
                    }),
            .out_data(lut_99_out)
        );

reg   lut_99_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_99_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_99_ff <= lut_99_out;
    end
end

assign out_data[99] = lut_99_ff;




// LUT : 100

wire lut_100_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100101101111100101110110111110111111000010101010111100111010),
            .DEVICE(DEVICE)
        )
    i_lut_100
        (
            .in_data({
                         in_data[74],
                         in_data[385],
                         in_data[562],
                         in_data[697],
                         in_data[357],
                         in_data[567]
                    }),
            .out_data(lut_100_out)
        );

reg   lut_100_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_100_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_100_ff <= lut_100_out;
    end
end

assign out_data[100] = lut_100_ff;




// LUT : 101

wire lut_101_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011111010110011010111010101010011110101101000110000010111100),
            .DEVICE(DEVICE)
        )
    i_lut_101
        (
            .in_data({
                         in_data[46],
                         in_data[103],
                         in_data[698],
                         in_data[135],
                         in_data[8],
                         in_data[621]
                    }),
            .out_data(lut_101_out)
        );

reg   lut_101_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_101_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_101_ff <= lut_101_out;
    end
end

assign out_data[101] = lut_101_ff;




// LUT : 102

wire lut_102_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010011111000110110100100100001000000101100010111010101010011),
            .DEVICE(DEVICE)
        )
    i_lut_102
        (
            .in_data({
                         in_data[541],
                         in_data[668],
                         in_data[641],
                         in_data[479],
                         in_data[769],
                         in_data[682]
                    }),
            .out_data(lut_102_out)
        );

reg   lut_102_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_102_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_102_ff <= lut_102_out;
    end
end

assign out_data[102] = lut_102_ff;




// LUT : 103

wire lut_103_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111011111111001000110000001100011001110001010000101101111110),
            .DEVICE(DEVICE)
        )
    i_lut_103
        (
            .in_data({
                         in_data[675],
                         in_data[618],
                         in_data[120],
                         in_data[588],
                         in_data[363],
                         in_data[447]
                    }),
            .out_data(lut_103_out)
        );

reg   lut_103_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_103_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_103_ff <= lut_103_out;
    end
end

assign out_data[103] = lut_103_ff;




// LUT : 104

wire lut_104_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001010000011101100000111010101000100010001000111011010000100),
            .DEVICE(DEVICE)
        )
    i_lut_104
        (
            .in_data({
                         in_data[235],
                         in_data[52],
                         in_data[411],
                         in_data[558],
                         in_data[287],
                         in_data[140]
                    }),
            .out_data(lut_104_out)
        );

reg   lut_104_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_104_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_104_ff <= lut_104_out;
    end
end

assign out_data[104] = lut_104_ff;




// LUT : 105

wire lut_105_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011100010001010011111001000101000011001100110110111110000011),
            .DEVICE(DEVICE)
        )
    i_lut_105
        (
            .in_data({
                         in_data[496],
                         in_data[244],
                         in_data[715],
                         in_data[553],
                         in_data[127],
                         in_data[194]
                    }),
            .out_data(lut_105_out)
        );

reg   lut_105_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_105_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_105_ff <= lut_105_out;
    end
end

assign out_data[105] = lut_105_ff;




// LUT : 106

wire lut_106_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100101111111001111101111110100111000100111101000111010011111),
            .DEVICE(DEVICE)
        )
    i_lut_106
        (
            .in_data({
                         in_data[515],
                         in_data[737],
                         in_data[636],
                         in_data[87],
                         in_data[227],
                         in_data[688]
                    }),
            .out_data(lut_106_out)
        );

reg   lut_106_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_106_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_106_ff <= lut_106_out;
    end
end

assign out_data[106] = lut_106_ff;




// LUT : 107

wire lut_107_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101011110101001100000101100011011010110011000110111000110011),
            .DEVICE(DEVICE)
        )
    i_lut_107
        (
            .in_data({
                         in_data[50],
                         in_data[768],
                         in_data[188],
                         in_data[498],
                         in_data[772],
                         in_data[240]
                    }),
            .out_data(lut_107_out)
        );

reg   lut_107_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_107_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_107_ff <= lut_107_out;
    end
end

assign out_data[107] = lut_107_ff;




// LUT : 108

wire lut_108_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111100101001100101111001101111110000011110000111001110010111111),
            .DEVICE(DEVICE)
        )
    i_lut_108
        (
            .in_data({
                         in_data[569],
                         in_data[716],
                         in_data[349],
                         in_data[476],
                         in_data[532],
                         in_data[202]
                    }),
            .out_data(lut_108_out)
        );

reg   lut_108_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_108_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_108_ff <= lut_108_out;
    end
end

assign out_data[108] = lut_108_ff;




// LUT : 109

wire lut_109_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101000001111101101011001001101100011000010011101001010110111),
            .DEVICE(DEVICE)
        )
    i_lut_109
        (
            .in_data({
                         in_data[722],
                         in_data[691],
                         in_data[556],
                         in_data[36],
                         in_data[72],
                         in_data[115]
                    }),
            .out_data(lut_109_out)
        );

reg   lut_109_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_109_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_109_ff <= lut_109_out;
    end
end

assign out_data[109] = lut_109_ff;




// LUT : 110

wire lut_110_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011010111111101111111111110111101000101111011001101011100101110),
            .DEVICE(DEVICE)
        )
    i_lut_110
        (
            .in_data({
                         in_data[469],
                         in_data[734],
                         in_data[133],
                         in_data[597],
                         in_data[438],
                         in_data[273]
                    }),
            .out_data(lut_110_out)
        );

reg   lut_110_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_110_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_110_ff <= lut_110_out;
    end
end

assign out_data[110] = lut_110_ff;




// LUT : 111

wire lut_111_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100011110111111110111100101010111011101011111011010001011100100),
            .DEVICE(DEVICE)
        )
    i_lut_111
        (
            .in_data({
                         in_data[308],
                         in_data[124],
                         in_data[259],
                         in_data[315],
                         in_data[430],
                         in_data[253]
                    }),
            .out_data(lut_111_out)
        );

reg   lut_111_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_111_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_111_ff <= lut_111_out;
    end
end

assign out_data[111] = lut_111_ff;




// LUT : 112

wire lut_112_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010110111100011011001011000000111111110011000111001110110110),
            .DEVICE(DEVICE)
        )
    i_lut_112
        (
            .in_data({
                         in_data[278],
                         in_data[660],
                         in_data[118],
                         in_data[121],
                         in_data[615],
                         in_data[90]
                    }),
            .out_data(lut_112_out)
        );

reg   lut_112_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_112_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_112_ff <= lut_112_out;
    end
end

assign out_data[112] = lut_112_ff;




// LUT : 113

wire lut_113_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100010010010111001111110011111111010110000010011000111010011010),
            .DEVICE(DEVICE)
        )
    i_lut_113
        (
            .in_data({
                         in_data[493],
                         in_data[85],
                         in_data[81],
                         in_data[282],
                         in_data[157],
                         in_data[80]
                    }),
            .out_data(lut_113_out)
        );

reg   lut_113_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_113_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_113_ff <= lut_113_out;
    end
end

assign out_data[113] = lut_113_ff;




// LUT : 114

wire lut_114_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101011101000010001110111100000000010010001110000111110101011),
            .DEVICE(DEVICE)
        )
    i_lut_114
        (
            .in_data({
                         in_data[224],
                         in_data[78],
                         in_data[248],
                         in_data[230],
                         in_data[654],
                         in_data[153]
                    }),
            .out_data(lut_114_out)
        );

reg   lut_114_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_114_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_114_ff <= lut_114_out;
    end
end

assign out_data[114] = lut_114_ff;




// LUT : 115

wire lut_115_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100101011011000110010111100110010011011110110100010011100100100),
            .DEVICE(DEVICE)
        )
    i_lut_115
        (
            .in_data({
                         in_data[198],
                         in_data[752],
                         in_data[258],
                         in_data[10],
                         in_data[761],
                         in_data[376]
                    }),
            .out_data(lut_115_out)
        );

reg   lut_115_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_115_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_115_ff <= lut_115_out;
    end
end

assign out_data[115] = lut_115_ff;




// LUT : 116

wire lut_116_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100101010101010010010011110010110110011001111000011000001110),
            .DEVICE(DEVICE)
        )
    i_lut_116
        (
            .in_data({
                         in_data[112],
                         in_data[27],
                         in_data[30],
                         in_data[559],
                         in_data[685],
                         in_data[275]
                    }),
            .out_data(lut_116_out)
        );

reg   lut_116_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_116_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_116_ff <= lut_116_out;
    end
end

assign out_data[116] = lut_116_ff;




// LUT : 117

wire lut_117_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100001110001100100000000000101000111110011110010010101011101),
            .DEVICE(DEVICE)
        )
    i_lut_117
        (
            .in_data({
                         in_data[546],
                         in_data[760],
                         in_data[550],
                         in_data[723],
                         in_data[594],
                         in_data[557]
                    }),
            .out_data(lut_117_out)
        );

reg   lut_117_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_117_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_117_ff <= lut_117_out;
    end
end

assign out_data[117] = lut_117_ff;




// LUT : 118

wire lut_118_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001011111011110000010111111000101101101010110011111010001110),
            .DEVICE(DEVICE)
        )
    i_lut_118
        (
            .in_data({
                         in_data[612],
                         in_data[542],
                         in_data[780],
                         in_data[274],
                         in_data[177],
                         in_data[182]
                    }),
            .out_data(lut_118_out)
        );

reg   lut_118_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_118_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_118_ff <= lut_118_out;
    end
end

assign out_data[118] = lut_118_ff;




// LUT : 119

wire lut_119_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000010010100001111000011100001001001101010010100100100000001),
            .DEVICE(DEVICE)
        )
    i_lut_119
        (
            .in_data({
                         in_data[645],
                         in_data[519],
                         in_data[412],
                         in_data[700],
                         in_data[285],
                         in_data[450]
                    }),
            .out_data(lut_119_out)
        );

reg   lut_119_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_119_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_119_ff <= lut_119_out;
    end
end

assign out_data[119] = lut_119_ff;




// LUT : 120

wire lut_120_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010111001101011111000010101011001101100011101100011110001000),
            .DEVICE(DEVICE)
        )
    i_lut_120
        (
            .in_data({
                         in_data[425],
                         in_data[241],
                         in_data[743],
                         in_data[205],
                         in_data[383],
                         in_data[9]
                    }),
            .out_data(lut_120_out)
        );

reg   lut_120_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_120_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_120_ff <= lut_120_out;
    end
end

assign out_data[120] = lut_120_ff;




// LUT : 121

wire lut_121_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000000100010100101111110111100111110111000110010100010010000),
            .DEVICE(DEVICE)
        )
    i_lut_121
        (
            .in_data({
                         in_data[644],
                         in_data[57],
                         in_data[38],
                         in_data[464],
                         in_data[676],
                         in_data[366]
                    }),
            .out_data(lut_121_out)
        );

reg   lut_121_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_121_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_121_ff <= lut_121_out;
    end
end

assign out_data[121] = lut_121_ff;




// LUT : 122

wire lut_122_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111101001001110001011101001000111110111000110010010000110101),
            .DEVICE(DEVICE)
        )
    i_lut_122
        (
            .in_data({
                         in_data[233],
                         in_data[643],
                         in_data[264],
                         in_data[503],
                         in_data[599],
                         in_data[748]
                    }),
            .out_data(lut_122_out)
        );

reg   lut_122_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_122_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_122_ff <= lut_122_out;
    end
end

assign out_data[122] = lut_122_ff;




// LUT : 123

wire lut_123_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000110011011100010111000111111110000011101110110111101001111110),
            .DEVICE(DEVICE)
        )
    i_lut_123
        (
            .in_data({
                         in_data[712],
                         in_data[669],
                         in_data[329],
                         in_data[199],
                         in_data[468],
                         in_data[708]
                    }),
            .out_data(lut_123_out)
        );

reg   lut_123_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_123_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_123_ff <= lut_123_out;
    end
end

assign out_data[123] = lut_123_ff;




// LUT : 124

wire lut_124_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110100111111100110110111011001000111101001001011111011101000),
            .DEVICE(DEVICE)
        )
    i_lut_124
        (
            .in_data({
                         in_data[319],
                         in_data[312],
                         in_data[145],
                         in_data[683],
                         in_data[477],
                         in_data[354]
                    }),
            .out_data(lut_124_out)
        );

reg   lut_124_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_124_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_124_ff <= lut_124_out;
    end
end

assign out_data[124] = lut_124_ff;




// LUT : 125

wire lut_125_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010001010111101011111010000101110001100100111011010001110011),
            .DEVICE(DEVICE)
        )
    i_lut_125
        (
            .in_data({
                         in_data[555],
                         in_data[344],
                         in_data[656],
                         in_data[747],
                         in_data[563],
                         in_data[250]
                    }),
            .out_data(lut_125_out)
        );

reg   lut_125_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_125_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_125_ff <= lut_125_out;
    end
end

assign out_data[125] = lut_125_ff;




// LUT : 126

wire lut_126_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110001100010010001101010001010110111000011001110010110001111),
            .DEVICE(DEVICE)
        )
    i_lut_126
        (
            .in_data({
                         in_data[47],
                         in_data[735],
                         in_data[661],
                         in_data[711],
                         in_data[24],
                         in_data[197]
                    }),
            .out_data(lut_126_out)
        );

reg   lut_126_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_126_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_126_ff <= lut_126_out;
    end
end

assign out_data[126] = lut_126_ff;




// LUT : 127

wire lut_127_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010001111001100000000001000011000100010100010101000000010000),
            .DEVICE(DEVICE)
        )
    i_lut_127
        (
            .in_data({
                         in_data[263],
                         in_data[159],
                         in_data[613],
                         in_data[48],
                         in_data[505],
                         in_data[625]
                    }),
            .out_data(lut_127_out)
        );

reg   lut_127_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_127_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_127_ff <= lut_127_out;
    end
end

assign out_data[127] = lut_127_ff;




// LUT : 128

wire lut_128_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000000110101001000001011100001000100000000001001000010000100),
            .DEVICE(DEVICE)
        )
    i_lut_128
        (
            .in_data({
                         in_data[34],
                         in_data[443],
                         in_data[525],
                         in_data[631],
                         in_data[407],
                         in_data[356]
                    }),
            .out_data(lut_128_out)
        );

reg   lut_128_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_128_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_128_ff <= lut_128_out;
    end
end

assign out_data[128] = lut_128_ff;




// LUT : 129

wire lut_129_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010010001110100110000001111010100100001001110001100011101000101),
            .DEVICE(DEVICE)
        )
    i_lut_129
        (
            .in_data({
                         in_data[189],
                         in_data[88],
                         in_data[348],
                         in_data[730],
                         in_data[517],
                         in_data[346]
                    }),
            .out_data(lut_129_out)
        );

reg   lut_129_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_129_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_129_ff <= lut_129_out;
    end
end

assign out_data[129] = lut_129_ff;




// LUT : 130

wire lut_130_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111111010111111101110111001100111101000011100111011100010010),
            .DEVICE(DEVICE)
        )
    i_lut_130
        (
            .in_data({
                         in_data[257],
                         in_data[433],
                         in_data[659],
                         in_data[16],
                         in_data[144],
                         in_data[766]
                    }),
            .out_data(lut_130_out)
        );

reg   lut_130_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_130_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_130_ff <= lut_130_out;
    end
end

assign out_data[130] = lut_130_ff;




// LUT : 131

wire lut_131_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111111100001001110101110111000011111011101011000111011101110),
            .DEVICE(DEVICE)
        )
    i_lut_131
        (
            .in_data({
                         in_data[417],
                         in_data[172],
                         in_data[689],
                         in_data[641],
                         in_data[410],
                         in_data[743]
                    }),
            .out_data(lut_131_out)
        );

reg   lut_131_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_131_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_131_ff <= lut_131_out;
    end
end

assign out_data[131] = lut_131_ff;




// LUT : 132

wire lut_132_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001101100010011010011000111001011010101001011011011100000110000),
            .DEVICE(DEVICE)
        )
    i_lut_132
        (
            .in_data({
                         in_data[32],
                         in_data[103],
                         in_data[521],
                         in_data[194],
                         in_data[419],
                         in_data[693]
                    }),
            .out_data(lut_132_out)
        );

reg   lut_132_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_132_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_132_ff <= lut_132_out;
    end
end

assign out_data[132] = lut_132_ff;




// LUT : 133

wire lut_133_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100000100000000000110001111010000000001001011000101110000110),
            .DEVICE(DEVICE)
        )
    i_lut_133
        (
            .in_data({
                         in_data[509],
                         in_data[129],
                         in_data[122],
                         in_data[649],
                         in_data[127],
                         in_data[82]
                    }),
            .out_data(lut_133_out)
        );

reg   lut_133_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_133_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_133_ff <= lut_133_out;
    end
end

assign out_data[133] = lut_133_ff;




// LUT : 134

wire lut_134_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111101000100110011110011101000000100010101010000100001011011),
            .DEVICE(DEVICE)
        )
    i_lut_134
        (
            .in_data({
                         in_data[552],
                         in_data[191],
                         in_data[101],
                         in_data[602],
                         in_data[578],
                         in_data[549]
                    }),
            .out_data(lut_134_out)
        );

reg   lut_134_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_134_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_134_ff <= lut_134_out;
    end
end

assign out_data[134] = lut_134_ff;




// LUT : 135

wire lut_135_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001000000010100010100111101011101111111111101111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_135
        (
            .in_data({
                         in_data[655],
                         in_data[604],
                         in_data[398],
                         in_data[405],
                         in_data[107],
                         in_data[454]
                    }),
            .out_data(lut_135_out)
        );

reg   lut_135_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_135_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_135_ff <= lut_135_out;
    end
end

assign out_data[135] = lut_135_ff;




// LUT : 136

wire lut_136_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100101000100001101000011101001111101111100000110110001100110011),
            .DEVICE(DEVICE)
        )
    i_lut_136
        (
            .in_data({
                         in_data[275],
                         in_data[138],
                         in_data[494],
                         in_data[363],
                         in_data[382],
                         in_data[514]
                    }),
            .out_data(lut_136_out)
        );

reg   lut_136_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_136_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_136_ff <= lut_136_out;
    end
end

assign out_data[136] = lut_136_ff;




// LUT : 137

wire lut_137_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111100101011101111111011101000001111011111110000011001110111),
            .DEVICE(DEVICE)
        )
    i_lut_137
        (
            .in_data({
                         in_data[350],
                         in_data[440],
                         in_data[446],
                         in_data[577],
                         in_data[355],
                         in_data[407]
                    }),
            .out_data(lut_137_out)
        );

reg   lut_137_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_137_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_137_ff <= lut_137_out;
    end
end

assign out_data[137] = lut_137_ff;




// LUT : 138

wire lut_138_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010111111101111010011110111111110111010010110100000101111011010),
            .DEVICE(DEVICE)
        )
    i_lut_138
        (
            .in_data({
                         in_data[348],
                         in_data[159],
                         in_data[330],
                         in_data[478],
                         in_data[187],
                         in_data[222]
                    }),
            .out_data(lut_138_out)
        );

reg   lut_138_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_138_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_138_ff <= lut_138_out;
    end
end

assign out_data[138] = lut_138_ff;




// LUT : 139

wire lut_139_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101101001101000101111010010001001111100001011011100100101100),
            .DEVICE(DEVICE)
        )
    i_lut_139
        (
            .in_data({
                         in_data[459],
                         in_data[169],
                         in_data[105],
                         in_data[346],
                         in_data[682],
                         in_data[111]
                    }),
            .out_data(lut_139_out)
        );

reg   lut_139_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_139_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_139_ff <= lut_139_out;
    end
end

assign out_data[139] = lut_139_ff;




// LUT : 140

wire lut_140_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011100111101100101101001011111100011001010001001000011010101),
            .DEVICE(DEVICE)
        )
    i_lut_140
        (
            .in_data({
                         in_data[125],
                         in_data[227],
                         in_data[43],
                         in_data[112],
                         in_data[722],
                         in_data[277]
                    }),
            .out_data(lut_140_out)
        );

reg   lut_140_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_140_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_140_ff <= lut_140_out;
    end
end

assign out_data[140] = lut_140_ff;




// LUT : 141

wire lut_141_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100010101011011001001110111111000001011111011011111011010101),
            .DEVICE(DEVICE)
        )
    i_lut_141
        (
            .in_data({
                         in_data[607],
                         in_data[550],
                         in_data[768],
                         in_data[268],
                         in_data[49],
                         in_data[751]
                    }),
            .out_data(lut_141_out)
        );

reg   lut_141_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_141_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_141_ff <= lut_141_out;
    end
end

assign out_data[141] = lut_141_ff;




// LUT : 142

wire lut_142_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110000110011011011001111111111100101101001100000100101001101),
            .DEVICE(DEVICE)
        )
    i_lut_142
        (
            .in_data({
                         in_data[210],
                         in_data[67],
                         in_data[51],
                         in_data[519],
                         in_data[628],
                         in_data[412]
                    }),
            .out_data(lut_142_out)
        );

reg   lut_142_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_142_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_142_ff <= lut_142_out;
    end
end

assign out_data[142] = lut_142_ff;




// LUT : 143

wire lut_143_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000110010000010111110110111000110000110101100101011111111110),
            .DEVICE(DEVICE)
        )
    i_lut_143
        (
            .in_data({
                         in_data[713],
                         in_data[143],
                         in_data[195],
                         in_data[538],
                         in_data[192],
                         in_data[276]
                    }),
            .out_data(lut_143_out)
        );

reg   lut_143_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_143_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_143_ff <= lut_143_out;
    end
end

assign out_data[143] = lut_143_ff;




// LUT : 144

wire lut_144_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001110011000111101111100110111111110011001000001011011110001001),
            .DEVICE(DEVICE)
        )
    i_lut_144
        (
            .in_data({
                         in_data[301],
                         in_data[531],
                         in_data[364],
                         in_data[124],
                         in_data[706],
                         in_data[623]
                    }),
            .out_data(lut_144_out)
        );

reg   lut_144_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_144_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_144_ff <= lut_144_out;
    end
end

assign out_data[144] = lut_144_ff;




// LUT : 145

wire lut_145_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011111000101001000101000010110111100101100010011101010000000),
            .DEVICE(DEVICE)
        )
    i_lut_145
        (
            .in_data({
                         in_data[597],
                         in_data[598],
                         in_data[36],
                         in_data[564],
                         in_data[240],
                         in_data[366]
                    }),
            .out_data(lut_145_out)
        );

reg   lut_145_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_145_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_145_ff <= lut_145_out;
    end
end

assign out_data[145] = lut_145_ff;




// LUT : 146

wire lut_146_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001111110101000100011011100100000001000000110101001000100001001),
            .DEVICE(DEVICE)
        )
    i_lut_146
        (
            .in_data({
                         in_data[500],
                         in_data[736],
                         in_data[344],
                         in_data[85],
                         in_data[735],
                         in_data[118]
                    }),
            .out_data(lut_146_out)
        );

reg   lut_146_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_146_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_146_ff <= lut_146_out;
    end
end

assign out_data[146] = lut_146_ff;




// LUT : 147

wire lut_147_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001010100111101110001111000110010001010100010000001111010111),
            .DEVICE(DEVICE)
        )
    i_lut_147
        (
            .in_data({
                         in_data[283],
                         in_data[90],
                         in_data[116],
                         in_data[753],
                         in_data[762],
                         in_data[698]
                    }),
            .out_data(lut_147_out)
        );

reg   lut_147_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_147_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_147_ff <= lut_147_out;
    end
end

assign out_data[147] = lut_147_ff;




// LUT : 148

wire lut_148_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101111110100101110111010110010010100010110100111010101101100),
            .DEVICE(DEVICE)
        )
    i_lut_148
        (
            .in_data({
                         in_data[428],
                         in_data[207],
                         in_data[445],
                         in_data[455],
                         in_data[477],
                         in_data[223]
                    }),
            .out_data(lut_148_out)
        );

reg   lut_148_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_148_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_148_ff <= lut_148_out;
    end
end

assign out_data[148] = lut_148_ff;




// LUT : 149

wire lut_149_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000101101111000000000000000000010000000100000010000011100000),
            .DEVICE(DEVICE)
        )
    i_lut_149
        (
            .in_data({
                         in_data[77],
                         in_data[763],
                         in_data[400],
                         in_data[525],
                         in_data[236],
                         in_data[465]
                    }),
            .out_data(lut_149_out)
        );

reg   lut_149_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_149_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_149_ff <= lut_149_out;
    end
end

assign out_data[149] = lut_149_ff;




// LUT : 150

wire lut_150_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000001110100111101011100110101110111111011001111111111001100),
            .DEVICE(DEVICE)
        )
    i_lut_150
        (
            .in_data({
                         in_data[453],
                         in_data[183],
                         in_data[594],
                         in_data[320],
                         in_data[100],
                         in_data[367]
                    }),
            .out_data(lut_150_out)
        );

reg   lut_150_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_150_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_150_ff <= lut_150_out;
    end
end

assign out_data[150] = lut_150_ff;




// LUT : 151

wire lut_151_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110110100010101011101001100101100011110111101110010100111011111),
            .DEVICE(DEVICE)
        )
    i_lut_151
        (
            .in_data({
                         in_data[390],
                         in_data[420],
                         in_data[12],
                         in_data[273],
                         in_data[337],
                         in_data[186]
                    }),
            .out_data(lut_151_out)
        );

reg   lut_151_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_151_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_151_ff <= lut_151_out;
    end
end

assign out_data[151] = lut_151_ff;




// LUT : 152

wire lut_152_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100001010110101011001001101000011110001011111001101100001111),
            .DEVICE(DEVICE)
        )
    i_lut_152
        (
            .in_data({
                         in_data[738],
                         in_data[451],
                         in_data[640],
                         in_data[74],
                         in_data[220],
                         in_data[136]
                    }),
            .out_data(lut_152_out)
        );

reg   lut_152_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_152_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_152_ff <= lut_152_out;
    end
end

assign out_data[152] = lut_152_ff;




// LUT : 153

wire lut_153_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101011111010000101100010011011010110110111110001011011010111),
            .DEVICE(DEVICE)
        )
    i_lut_153
        (
            .in_data({
                         in_data[461],
                         in_data[151],
                         in_data[485],
                         in_data[165],
                         in_data[721],
                         in_data[254]
                    }),
            .out_data(lut_153_out)
        );

reg   lut_153_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_153_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_153_ff <= lut_153_out;
    end
end

assign out_data[153] = lut_153_ff;




// LUT : 154

wire lut_154_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111111110111011101111111010101010100100),
            .DEVICE(DEVICE)
        )
    i_lut_154
        (
            .in_data({
                         in_data[584],
                         in_data[260],
                         in_data[324],
                         in_data[299],
                         in_data[234],
                         in_data[583]
                    }),
            .out_data(lut_154_out)
        );

reg   lut_154_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_154_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_154_ff <= lut_154_out;
    end
end

assign out_data[154] = lut_154_ff;




// LUT : 155

wire lut_155_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111101010010000010000100010001110110011101101000010010100101),
            .DEVICE(DEVICE)
        )
    i_lut_155
        (
            .in_data({
                         in_data[650],
                         in_data[18],
                         in_data[131],
                         in_data[161],
                         in_data[671],
                         in_data[319]
                    }),
            .out_data(lut_155_out)
        );

reg   lut_155_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_155_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_155_ff <= lut_155_out;
    end
end

assign out_data[155] = lut_155_ff;




// LUT : 156

wire lut_156_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001111101010101111001011010010101010000101001001010010010100),
            .DEVICE(DEVICE)
        )
    i_lut_156
        (
            .in_data({
                         in_data[486],
                         in_data[25],
                         in_data[188],
                         in_data[84],
                         in_data[632],
                         in_data[568]
                    }),
            .out_data(lut_156_out)
        );

reg   lut_156_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_156_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_156_ff <= lut_156_out;
    end
end

assign out_data[156] = lut_156_ff;




// LUT : 157

wire lut_157_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000110110011011111001111000101111111001100011011011110110001),
            .DEVICE(DEVICE)
        )
    i_lut_157
        (
            .in_data({
                         in_data[378],
                         in_data[269],
                         in_data[388],
                         in_data[360],
                         in_data[696],
                         in_data[467]
                    }),
            .out_data(lut_157_out)
        );

reg   lut_157_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_157_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_157_ff <= lut_157_out;
    end
end

assign out_data[157] = lut_157_ff;




// LUT : 158

wire lut_158_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111100000100001101111011001100011000111111011001101100110011),
            .DEVICE(DEVICE)
        )
    i_lut_158
        (
            .in_data({
                         in_data[300],
                         in_data[8],
                         in_data[776],
                         in_data[289],
                         in_data[387],
                         in_data[562]
                    }),
            .out_data(lut_158_out)
        );

reg   lut_158_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_158_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_158_ff <= lut_158_out;
    end
end

assign out_data[158] = lut_158_ff;




// LUT : 159

wire lut_159_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001011001111101101001100110001001100011010001101010001110100),
            .DEVICE(DEVICE)
        )
    i_lut_159
        (
            .in_data({
                         in_data[152],
                         in_data[23],
                         in_data[353],
                         in_data[755],
                         in_data[517],
                         in_data[57]
                    }),
            .out_data(lut_159_out)
        );

reg   lut_159_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_159_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_159_ff <= lut_159_out;
    end
end

assign out_data[159] = lut_159_ff;




// LUT : 160

wire lut_160_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010110001000000000001000100111111111100011100001101001101000111),
            .DEVICE(DEVICE)
        )
    i_lut_160
        (
            .in_data({
                         in_data[690],
                         in_data[371],
                         in_data[427],
                         in_data[647],
                         in_data[560],
                         in_data[380]
                    }),
            .out_data(lut_160_out)
        );

reg   lut_160_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_160_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_160_ff <= lut_160_out;
    end
end

assign out_data[160] = lut_160_ff;




// LUT : 161

wire lut_161_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110111110000010111100011101011011000000010001000110010011111110),
            .DEVICE(DEVICE)
        )
    i_lut_161
        (
            .in_data({
                         in_data[757],
                         in_data[600],
                         in_data[312],
                         in_data[396],
                         in_data[190],
                         in_data[694]
                    }),
            .out_data(lut_161_out)
        );

reg   lut_161_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_161_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_161_ff <= lut_161_out;
    end
end

assign out_data[161] = lut_161_ff;




// LUT : 162

wire lut_162_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001001101001001001101101111110010000110011111110001100110011),
            .DEVICE(DEVICE)
        )
    i_lut_162
        (
            .in_data({
                         in_data[644],
                         in_data[677],
                         in_data[544],
                         in_data[339],
                         in_data[401],
                         in_data[354]
                    }),
            .out_data(lut_162_out)
        );

reg   lut_162_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_162_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_162_ff <= lut_162_out;
    end
end

assign out_data[162] = lut_162_ff;




// LUT : 163

wire lut_163_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010010111011100110000001000100010100110101010011100000101001001),
            .DEVICE(DEVICE)
        )
    i_lut_163
        (
            .in_data({
                         in_data[466],
                         in_data[711],
                         in_data[158],
                         in_data[150],
                         in_data[45],
                         in_data[553]
                    }),
            .out_data(lut_163_out)
        );

reg   lut_163_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_163_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_163_ff <= lut_163_out;
    end
end

assign out_data[163] = lut_163_ff;




// LUT : 164

wire lut_164_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001011100100011000101110111000101010100011001110001110101011),
            .DEVICE(DEVICE)
        )
    i_lut_164
        (
            .in_data({
                         in_data[94],
                         in_data[515],
                         in_data[452],
                         in_data[267],
                         in_data[619],
                         in_data[29]
                    }),
            .out_data(lut_164_out)
        );

reg   lut_164_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_164_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_164_ff <= lut_164_out;
    end
end

assign out_data[164] = lut_164_ff;




// LUT : 165

wire lut_165_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001110101101010011010100110100110101011010110100110101001101),
            .DEVICE(DEVICE)
        )
    i_lut_165
        (
            .in_data({
                         in_data[237],
                         in_data[416],
                         in_data[574],
                         in_data[239],
                         in_data[590],
                         in_data[221]
                    }),
            .out_data(lut_165_out)
        );

reg   lut_165_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_165_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_165_ff <= lut_165_out;
    end
end

assign out_data[165] = lut_165_ff;




// LUT : 166

wire lut_166_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100010100000110011011000101010100101111011111010111100111011),
            .DEVICE(DEVICE)
        )
    i_lut_166
        (
            .in_data({
                         in_data[64],
                         in_data[464],
                         in_data[617],
                         in_data[147],
                         in_data[432],
                         in_data[679]
                    }),
            .out_data(lut_166_out)
        );

reg   lut_166_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_166_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_166_ff <= lut_166_out;
    end
end

assign out_data[166] = lut_166_ff;




// LUT : 167

wire lut_167_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100001101011110011101111111100000000001110001000110111110011),
            .DEVICE(DEVICE)
        )
    i_lut_167
        (
            .in_data({
                         in_data[724],
                         in_data[572],
                         in_data[153],
                         in_data[285],
                         in_data[206],
                         in_data[471]
                    }),
            .out_data(lut_167_out)
        );

reg   lut_167_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_167_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_167_ff <= lut_167_out;
    end
end

assign out_data[167] = lut_167_ff;




// LUT : 168

wire lut_168_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011010011111011110110010110100000111111111010110101110110101110),
            .DEVICE(DEVICE)
        )
    i_lut_168
        (
            .in_data({
                         in_data[727],
                         in_data[114],
                         in_data[702],
                         in_data[386],
                         in_data[712],
                         in_data[744]
                    }),
            .out_data(lut_168_out)
        );

reg   lut_168_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_168_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_168_ff <= lut_168_out;
    end
end

assign out_data[168] = lut_168_ff;




// LUT : 169

wire lut_169_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101010110010110111000110010001000010111100010110011100011000),
            .DEVICE(DEVICE)
        )
    i_lut_169
        (
            .in_data({
                         in_data[27],
                         in_data[566],
                         in_data[309],
                         in_data[139],
                         in_data[506],
                         in_data[444]
                    }),
            .out_data(lut_169_out)
        );

reg   lut_169_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_169_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_169_ff <= lut_169_out;
    end
end

assign out_data[169] = lut_169_ff;




// LUT : 170

wire lut_170_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001001011001110100001110110001101011100011111000000011111000),
            .DEVICE(DEVICE)
        )
    i_lut_170
        (
            .in_data({
                         in_data[493],
                         in_data[771],
                         in_data[304],
                         in_data[536],
                         in_data[245],
                         in_data[545]
                    }),
            .out_data(lut_170_out)
        );

reg   lut_170_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_170_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_170_ff <= lut_170_out;
    end
end

assign out_data[170] = lut_170_ff;




// LUT : 171

wire lut_171_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000001100111011010101100110000101010010100100000100011001111),
            .DEVICE(DEVICE)
        )
    i_lut_171
        (
            .in_data({
                         in_data[764],
                         in_data[55],
                         in_data[695],
                         in_data[662],
                         in_data[646],
                         in_data[342]
                    }),
            .out_data(lut_171_out)
        );

reg   lut_171_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_171_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_171_ff <= lut_171_out;
    end
end

assign out_data[171] = lut_171_ff;




// LUT : 172

wire lut_172_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001100001111010000011110100101100111000010010101010011111111111),
            .DEVICE(DEVICE)
        )
    i_lut_172
        (
            .in_data({
                         in_data[576],
                         in_data[97],
                         in_data[208],
                         in_data[672],
                         in_data[608],
                         in_data[133]
                    }),
            .out_data(lut_172_out)
        );

reg   lut_172_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_172_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_172_ff <= lut_172_out;
    end
end

assign out_data[172] = lut_172_ff;




// LUT : 173

wire lut_173_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010111000110010111101011101100010111010100110110101010110100),
            .DEVICE(DEVICE)
        )
    i_lut_173
        (
            .in_data({
                         in_data[431],
                         in_data[88],
                         in_data[703],
                         in_data[93],
                         in_data[612],
                         in_data[219]
                    }),
            .out_data(lut_173_out)
        );

reg   lut_173_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_173_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_173_ff <= lut_173_out;
    end
end

assign out_data[173] = lut_173_ff;




// LUT : 174

wire lut_174_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100101110111100100110101111101111101010001001001110101000101),
            .DEVICE(DEVICE)
        )
    i_lut_174
        (
            .in_data({
                         in_data[434],
                         in_data[154],
                         in_data[137],
                         in_data[331],
                         in_data[306],
                         in_data[481]
                    }),
            .out_data(lut_174_out)
        );

reg   lut_174_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_174_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_174_ff <= lut_174_out;
    end
end

assign out_data[174] = lut_174_ff;




// LUT : 175

wire lut_175_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000000100010011011010101101011000101101110110000100111000000),
            .DEVICE(DEVICE)
        )
    i_lut_175
        (
            .in_data({
                         in_data[228],
                         in_data[415],
                         in_data[395],
                         in_data[516],
                         in_data[266],
                         in_data[653]
                    }),
            .out_data(lut_175_out)
        );

reg   lut_175_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_175_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_175_ff <= lut_175_out;
    end
end

assign out_data[175] = lut_175_ff;




// LUT : 176

wire lut_176_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001011010110110111101011000011000111001110001010010111010000),
            .DEVICE(DEVICE)
        )
    i_lut_176
        (
            .in_data({
                         in_data[79],
                         in_data[134],
                         in_data[535],
                         in_data[7],
                         in_data[59],
                         in_data[687]
                    }),
            .out_data(lut_176_out)
        );

reg   lut_176_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_176_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_176_ff <= lut_176_out;
    end
end

assign out_data[176] = lut_176_ff;




// LUT : 177

wire lut_177_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111111101000000011110000100111011101010111111111000111110010),
            .DEVICE(DEVICE)
        )
    i_lut_177
        (
            .in_data({
                         in_data[274],
                         in_data[534],
                         in_data[651],
                         in_data[294],
                         in_data[205],
                         in_data[120]
                    }),
            .out_data(lut_177_out)
        );

reg   lut_177_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_177_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_177_ff <= lut_177_out;
    end
end

assign out_data[177] = lut_177_ff;




// LUT : 178

wire lut_178_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101111101110010111010110111011110001101010101010111011101110),
            .DEVICE(DEVICE)
        )
    i_lut_178
        (
            .in_data({
                         in_data[593],
                         in_data[209],
                         in_data[50],
                         in_data[264],
                         in_data[175],
                         in_data[462]
                    }),
            .out_data(lut_178_out)
        );

reg   lut_178_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_178_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_178_ff <= lut_178_out;
    end
end

assign out_data[178] = lut_178_ff;




// LUT : 179

wire lut_179_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010010100011001101000010000111111111001110010011100000000011101),
            .DEVICE(DEVICE)
        )
    i_lut_179
        (
            .in_data({
                         in_data[372],
                         in_data[335],
                         in_data[501],
                         in_data[758],
                         in_data[626],
                         in_data[463]
                    }),
            .out_data(lut_179_out)
        );

reg   lut_179_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_179_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_179_ff <= lut_179_out;
    end
end

assign out_data[179] = lut_179_ff;




// LUT : 180

wire lut_180_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010000101000110000000010010110001110000011000111111110001101),
            .DEVICE(DEVICE)
        )
    i_lut_180
        (
            .in_data({
                         in_data[760],
                         in_data[326],
                         in_data[162],
                         in_data[216],
                         in_data[767],
                         in_data[393]
                    }),
            .out_data(lut_180_out)
        );

reg   lut_180_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_180_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_180_ff <= lut_180_out;
    end
end

assign out_data[180] = lut_180_ff;




// LUT : 181

wire lut_181_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010100100111111101011100110010111000111100001010000101100000),
            .DEVICE(DEVICE)
        )
    i_lut_181
        (
            .in_data({
                         in_data[19],
                         in_data[730],
                         in_data[213],
                         in_data[476],
                         in_data[606],
                         in_data[76]
                    }),
            .out_data(lut_181_out)
        );

reg   lut_181_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_181_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_181_ff <= lut_181_out;
    end
end

assign out_data[181] = lut_181_ff;




// LUT : 182

wire lut_182_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011111100111111011010100011111010111010011110110000001010100),
            .DEVICE(DEVICE)
        )
    i_lut_182
        (
            .in_data({
                         in_data[773],
                         in_data[316],
                         in_data[343],
                         in_data[614],
                         in_data[265],
                         in_data[561]
                    }),
            .out_data(lut_182_out)
        );

reg   lut_182_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_182_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_182_ff <= lut_182_out;
    end
end

assign out_data[182] = lut_182_ff;




// LUT : 183

wire lut_183_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000000000000010000100000110011001000000011001110100000001100),
            .DEVICE(DEVICE)
        )
    i_lut_183
        (
            .in_data({
                         in_data[297],
                         in_data[551],
                         in_data[253],
                         in_data[480],
                         in_data[375],
                         in_data[149]
                    }),
            .out_data(lut_183_out)
        );

reg   lut_183_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_183_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_183_ff <= lut_183_out;
    end
end

assign out_data[183] = lut_183_ff;




// LUT : 184

wire lut_184_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000010110001011000100100001011100011110011010011111110101011),
            .DEVICE(DEVICE)
        )
    i_lut_184
        (
            .in_data({
                         in_data[504],
                         in_data[648],
                         in_data[484],
                         in_data[376],
                         in_data[505],
                         in_data[457]
                    }),
            .out_data(lut_184_out)
        );

reg   lut_184_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_184_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_184_ff <= lut_184_out;
    end
end

assign out_data[184] = lut_184_ff;




// LUT : 185

wire lut_185_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010011100111111110111011111011100100000101100100011111011111100),
            .DEVICE(DEVICE)
        )
    i_lut_185
        (
            .in_data({
                         in_data[66],
                         in_data[527],
                         in_data[352],
                         in_data[700],
                         in_data[414],
                         in_data[587]
                    }),
            .out_data(lut_185_out)
        );

reg   lut_185_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_185_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_185_ff <= lut_185_out;
    end
end

assign out_data[185] = lut_185_ff;




// LUT : 186

wire lut_186_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000110011010100110110010101101001000100010100101011000101011),
            .DEVICE(DEVICE)
        )
    i_lut_186
        (
            .in_data({
                         in_data[40],
                         in_data[745],
                         in_data[585],
                         in_data[307],
                         in_data[141],
                         in_data[438]
                    }),
            .out_data(lut_186_out)
        );

reg   lut_186_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_186_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_186_ff <= lut_186_out;
    end
end

assign out_data[186] = lut_186_ff;




// LUT : 187

wire lut_187_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101000000010000011010001100100011001101101111001101101111000),
            .DEVICE(DEVICE)
        )
    i_lut_187
        (
            .in_data({
                         in_data[252],
                         in_data[75],
                         in_data[557],
                         in_data[479],
                         in_data[196],
                         in_data[52]
                    }),
            .out_data(lut_187_out)
        );

reg   lut_187_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_187_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_187_ff <= lut_187_out;
    end
end

assign out_data[187] = lut_187_ff;




// LUT : 188

wire lut_188_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101111111010001110101001010101110101001100110100000010010001),
            .DEVICE(DEVICE)
        )
    i_lut_188
        (
            .in_data({
                         in_data[166],
                         in_data[176],
                         in_data[765],
                         in_data[513],
                         in_data[613],
                         in_data[365]
                    }),
            .out_data(lut_188_out)
        );

reg   lut_188_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_188_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_188_ff <= lut_188_out;
    end
end

assign out_data[188] = lut_188_ff;




// LUT : 189

wire lut_189_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000010111011011111111011111111111111010010001011001111011011),
            .DEVICE(DEVICE)
        )
    i_lut_189
        (
            .in_data({
                         in_data[171],
                         in_data[261],
                         in_data[63],
                         in_data[547],
                         in_data[756],
                         in_data[413]
                    }),
            .out_data(lut_189_out)
        );

reg   lut_189_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_189_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_189_ff <= lut_189_out;
    end
end

assign out_data[189] = lut_189_ff;




// LUT : 190

wire lut_190_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010011011100011010110000000010111001111111100110111000001001111),
            .DEVICE(DEVICE)
        )
    i_lut_190
        (
            .in_data({
                         in_data[246],
                         in_data[656],
                         in_data[9],
                         in_data[769],
                         in_data[759],
                         in_data[439]
                    }),
            .out_data(lut_190_out)
        );

reg   lut_190_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_190_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_190_ff <= lut_190_out;
    end
end

assign out_data[190] = lut_190_ff;




// LUT : 191

wire lut_191_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011011010101110001100110010011111010010000100000100101111011),
            .DEVICE(DEVICE)
        )
    i_lut_191
        (
            .in_data({
                         in_data[119],
                         in_data[35],
                         in_data[290],
                         in_data[115],
                         in_data[197],
                         in_data[422]
                    }),
            .out_data(lut_191_out)
        );

reg   lut_191_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_191_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_191_ff <= lut_191_out;
    end
end

assign out_data[191] = lut_191_ff;




// LUT : 192

wire lut_192_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000000110100000111001100011011001101100001010110100101101101),
            .DEVICE(DEVICE)
        )
    i_lut_192
        (
            .in_data({
                         in_data[603],
                         in_data[383],
                         in_data[146],
                         in_data[615],
                         in_data[775],
                         in_data[660]
                    }),
            .out_data(lut_192_out)
        );

reg   lut_192_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_192_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_192_ff <= lut_192_out;
    end
end

assign out_data[192] = lut_192_ff;




// LUT : 193

wire lut_193_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001000011110011101001111011100000111111101000110000100000101),
            .DEVICE(DEVICE)
        )
    i_lut_193
        (
            .in_data({
                         in_data[24],
                         in_data[643],
                         in_data[262],
                         in_data[750],
                         in_data[89],
                         in_data[739]
                    }),
            .out_data(lut_193_out)
        );

reg   lut_193_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_193_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_193_ff <= lut_193_out;
    end
end

assign out_data[193] = lut_193_ff;




// LUT : 194

wire lut_194_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110100001010111111010010011111111111101000100101010100100001),
            .DEVICE(DEVICE)
        )
    i_lut_194
        (
            .in_data({
                         in_data[621],
                         in_data[126],
                         in_data[323],
                         in_data[567],
                         in_data[148],
                         in_data[697]
                    }),
            .out_data(lut_194_out)
        );

reg   lut_194_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_194_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_194_ff <= lut_194_out;
    end
end

assign out_data[194] = lut_194_ff;




// LUT : 195

wire lut_195_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000100100010110110001010101110111110101110010001001010001101100),
            .DEVICE(DEVICE)
        )
    i_lut_195
        (
            .in_data({
                         in_data[22],
                         in_data[53],
                         in_data[540],
                         in_data[81],
                         in_data[20],
                         in_data[683]
                    }),
            .out_data(lut_195_out)
        );

reg   lut_195_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_195_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_195_ff <= lut_195_out;
    end
end

assign out_data[195] = lut_195_ff;




// LUT : 196

wire lut_196_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101001010001101110000010101111001101011101010101000011001000),
            .DEVICE(DEVICE)
        )
    i_lut_196
        (
            .in_data({
                         in_data[473],
                         in_data[322],
                         in_data[314],
                         in_data[46],
                         in_data[634],
                         in_data[3]
                    }),
            .out_data(lut_196_out)
        );

reg   lut_196_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_196_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_196_ff <= lut_196_out;
    end
end

assign out_data[196] = lut_196_ff;




// LUT : 197

wire lut_197_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110100000000000100000000000000101000000001010000010010000101),
            .DEVICE(DEVICE)
        )
    i_lut_197
        (
            .in_data({
                         in_data[498],
                         in_data[332],
                         in_data[620],
                         in_data[179],
                         in_data[347],
                         in_data[385]
                    }),
            .out_data(lut_197_out)
        );

reg   lut_197_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_197_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_197_ff <= lut_197_out;
    end
end

assign out_data[197] = lut_197_ff;




// LUT : 198

wire lut_198_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011011100101100001111110010110001101011001100000001110110101100),
            .DEVICE(DEVICE)
        )
    i_lut_198
        (
            .in_data({
                         in_data[145],
                         in_data[255],
                         in_data[408],
                         in_data[113],
                         in_data[315],
                         in_data[539]
                    }),
            .out_data(lut_198_out)
        );

reg   lut_198_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_198_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_198_ff <= lut_198_out;
    end
end

assign out_data[198] = lut_198_ff;




// LUT : 199

wire lut_199_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000010111111010100110101111111111111111111111101111111010000),
            .DEVICE(DEVICE)
        )
    i_lut_199
        (
            .in_data({
                         in_data[70],
                         in_data[573],
                         in_data[303],
                         in_data[678],
                         in_data[204],
                         in_data[328]
                    }),
            .out_data(lut_199_out)
        );

reg   lut_199_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_199_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_199_ff <= lut_199_out;
    end
end

assign out_data[199] = lut_199_ff;




// LUT : 200

wire lut_200_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001001011010111100111111011101000110110110110100011000110),
            .DEVICE(DEVICE)
        )
    i_lut_200
        (
            .in_data({
                         in_data[44],
                         in_data[726],
                         in_data[167],
                         in_data[708],
                         in_data[605],
                         in_data[394]
                    }),
            .out_data(lut_200_out)
        );

reg   lut_200_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_200_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_200_ff <= lut_200_out;
    end
end

assign out_data[200] = lut_200_ff;




// LUT : 201

wire lut_201_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000111100010010110010010000011110100100110011110000010100101),
            .DEVICE(DEVICE)
        )
    i_lut_201
        (
            .in_data({
                         in_data[110],
                         in_data[281],
                         in_data[748],
                         in_data[42],
                         in_data[201],
                         in_data[674]
                    }),
            .out_data(lut_201_out)
        );

reg   lut_201_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_201_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_201_ff <= lut_201_out;
    end
end

assign out_data[201] = lut_201_ff;




// LUT : 202

wire lut_202_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100011100010111110000110101110111111111111101111111100001100),
            .DEVICE(DEVICE)
        )
    i_lut_202
        (
            .in_data({
                         in_data[135],
                         in_data[482],
                         in_data[123],
                         in_data[520],
                         in_data[524],
                         in_data[259]
                    }),
            .out_data(lut_202_out)
        );

reg   lut_202_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_202_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_202_ff <= lut_202_out;
    end
end

assign out_data[202] = lut_202_ff;




// LUT : 203

wire lut_203_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110100001110110011101110111000000001001001011110110111101011),
            .DEVICE(DEVICE)
        )
    i_lut_203
        (
            .in_data({
                         in_data[178],
                         in_data[533],
                         in_data[510],
                         in_data[241],
                         in_data[443],
                         in_data[218]
                    }),
            .out_data(lut_203_out)
        );

reg   lut_203_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_203_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_203_ff <= lut_203_out;
    end
end

assign out_data[203] = lut_203_ff;




// LUT : 204

wire lut_204_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100111010100011100100110111111101111000001100111011011111100000),
            .DEVICE(DEVICE)
        )
    i_lut_204
        (
            .in_data({
                         in_data[117],
                         in_data[98],
                         in_data[1],
                         in_data[460],
                         in_data[507],
                         in_data[349]
                    }),
            .out_data(lut_204_out)
        );

reg   lut_204_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_204_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_204_ff <= lut_204_out;
    end
end

assign out_data[204] = lut_204_ff;




// LUT : 205

wire lut_205_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001001111100101111110101011001011101010110111111100000011001100),
            .DEVICE(DEVICE)
        )
    i_lut_205
        (
            .in_data({
                         in_data[142],
                         in_data[302],
                         in_data[174],
                         in_data[667],
                         in_data[272],
                         in_data[638]
                    }),
            .out_data(lut_205_out)
        );

reg   lut_205_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_205_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_205_ff <= lut_205_out;
    end
end

assign out_data[205] = lut_205_ff;




// LUT : 206

wire lut_206_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000010010110010111011111100101010001001111101000011110100000),
            .DEVICE(DEVICE)
        )
    i_lut_206
        (
            .in_data({
                         in_data[226],
                         in_data[670],
                         in_data[327],
                         in_data[95],
                         in_data[686],
                         in_data[106]
                    }),
            .out_data(lut_206_out)
        );

reg   lut_206_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_206_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_206_ff <= lut_206_out;
    end
end

assign out_data[206] = lut_206_ff;




// LUT : 207

wire lut_207_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110011001010111101001010111010011001010111011000100010000000),
            .DEVICE(DEVICE)
        )
    i_lut_207
        (
            .in_data({
                         in_data[778],
                         in_data[321],
                         in_data[406],
                         in_data[488],
                         in_data[503],
                         in_data[78]
                    }),
            .out_data(lut_207_out)
        );

reg   lut_207_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_207_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_207_ff <= lut_207_out;
    end
end

assign out_data[207] = lut_207_ff;




// LUT : 208

wire lut_208_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100111000101111010111110001011100101110010001010111111010101011),
            .DEVICE(DEVICE)
        )
    i_lut_208
        (
            .in_data({
                         in_data[173],
                         in_data[496],
                         in_data[546],
                         in_data[305],
                         in_data[10],
                         in_data[716]
                    }),
            .out_data(lut_208_out)
        );

reg   lut_208_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_208_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_208_ff <= lut_208_out;
    end
end

assign out_data[208] = lut_208_ff;




// LUT : 209

wire lut_209_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001101101101011011011111100101000101000011101011111111110000),
            .DEVICE(DEVICE)
        )
    i_lut_209
        (
            .in_data({
                         in_data[442],
                         in_data[637],
                         in_data[747],
                         in_data[68],
                         in_data[359],
                         in_data[155]
                    }),
            .out_data(lut_209_out)
        );

reg   lut_209_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_209_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_209_ff <= lut_209_out;
    end
end

assign out_data[209] = lut_209_ff;




// LUT : 210

wire lut_210_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100011000110011110001000111010000001010011111110100100011011),
            .DEVICE(DEVICE)
        )
    i_lut_210
        (
            .in_data({
                         in_data[13],
                         in_data[652],
                         in_data[15],
                         in_data[497],
                         in_data[73],
                         in_data[625]
                    }),
            .out_data(lut_210_out)
        );

reg   lut_210_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_210_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_210_ff <= lut_210_out;
    end
end

assign out_data[210] = lut_210_ff;




// LUT : 211

wire lut_211_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111000010100110011101110111010001000111111111100111011101110),
            .DEVICE(DEVICE)
        )
    i_lut_211
        (
            .in_data({
                         in_data[373],
                         in_data[170],
                         in_data[624],
                         in_data[468],
                         in_data[329],
                         in_data[357]
                    }),
            .out_data(lut_211_out)
        );

reg   lut_211_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_211_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_211_ff <= lut_211_out;
    end
end

assign out_data[211] = lut_211_ff;




// LUT : 212

wire lut_212_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010001111110010100010011110100111111110000100000100010010101),
            .DEVICE(DEVICE)
        )
    i_lut_212
        (
            .in_data({
                         in_data[421],
                         in_data[224],
                         in_data[458],
                         in_data[230],
                         in_data[308],
                         in_data[58]
                    }),
            .out_data(lut_212_out)
        );

reg   lut_212_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_212_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_212_ff <= lut_212_out;
    end
end

assign out_data[212] = lut_212_ff;




// LUT : 213

wire lut_213_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110110100000011110011011100000000110110110000011010010011110011),
            .DEVICE(DEVICE)
        )
    i_lut_213
        (
            .in_data({
                         in_data[669],
                         in_data[436],
                         in_data[774],
                         in_data[30],
                         in_data[668],
                         in_data[26]
                    }),
            .out_data(lut_213_out)
        );

reg   lut_213_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_213_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_213_ff <= lut_213_out;
    end
end

assign out_data[213] = lut_213_ff;




// LUT : 214

wire lut_214_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000110011111110001001011011111110111100000110001011100001011),
            .DEVICE(DEVICE)
        )
    i_lut_214
        (
            .in_data({
                         in_data[725],
                         in_data[180],
                         in_data[592],
                         in_data[489],
                         in_data[65],
                         in_data[635]
                    }),
            .out_data(lut_214_out)
        );

reg   lut_214_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_214_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_214_ff <= lut_214_out;
    end
end

assign out_data[214] = lut_214_ff;




// LUT : 215

wire lut_215_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100010100000011011000000111011000100010010110110000100001101),
            .DEVICE(DEVICE)
        )
    i_lut_215
        (
            .in_data({
                         in_data[714],
                         in_data[229],
                         in_data[636],
                         in_data[718],
                         in_data[588],
                         in_data[589]
                    }),
            .out_data(lut_215_out)
        );

reg   lut_215_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_215_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_215_ff <= lut_215_out;
    end
end

assign out_data[215] = lut_215_ff;




// LUT : 216

wire lut_216_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100010111100100101001011101011101001111111100000000110101000),
            .DEVICE(DEVICE)
        )
    i_lut_216
        (
            .in_data({
                         in_data[244],
                         in_data[313],
                         in_data[336],
                         in_data[379],
                         in_data[325],
                         in_data[742]
                    }),
            .out_data(lut_216_out)
        );

reg   lut_216_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_216_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_216_ff <= lut_216_out;
    end
end

assign out_data[216] = lut_216_ff;




// LUT : 217

wire lut_217_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000010001011110110101111101100001011110011111111101010111111),
            .DEVICE(DEVICE)
        )
    i_lut_217
        (
            .in_data({
                         in_data[580],
                         in_data[399],
                         in_data[542],
                         in_data[475],
                         in_data[575],
                         in_data[163]
                    }),
            .out_data(lut_217_out)
        );

reg   lut_217_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_217_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_217_ff <= lut_217_out;
    end
end

assign out_data[217] = lut_217_ff;




// LUT : 218

wire lut_218_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110100100011010100010110011011001000001000101111011010100010),
            .DEVICE(DEVICE)
        )
    i_lut_218
        (
            .in_data({
                         in_data[618],
                         in_data[160],
                         in_data[80],
                         in_data[263],
                         in_data[341],
                         in_data[491]
                    }),
            .out_data(lut_218_out)
        );

reg   lut_218_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_218_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_218_ff <= lut_218_out;
    end
end

assign out_data[218] = lut_218_ff;




// LUT : 219

wire lut_219_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010011111000000011110010110001101010111111010101010101100101011),
            .DEVICE(DEVICE)
        )
    i_lut_219
        (
            .in_data({
                         in_data[570],
                         in_data[291],
                         in_data[554],
                         in_data[38],
                         in_data[779],
                         in_data[0]
                    }),
            .out_data(lut_219_out)
        );

reg   lut_219_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_219_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_219_ff <= lut_219_out;
    end
end

assign out_data[219] = lut_219_ff;




// LUT : 220

wire lut_220_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001001100000010100001000110000000101111101011001010111110101110),
            .DEVICE(DEVICE)
        )
    i_lut_220
        (
            .in_data({
                         in_data[402],
                         in_data[437],
                         in_data[121],
                         in_data[391],
                         in_data[555],
                         in_data[599]
                    }),
            .out_data(lut_220_out)
        );

reg   lut_220_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_220_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_220_ff <= lut_220_out;
    end
end

assign out_data[220] = lut_220_ff;




// LUT : 221

wire lut_221_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100011000110111000001000100011010100010011111011000110011000011),
            .DEVICE(DEVICE)
        )
    i_lut_221
        (
            .in_data({
                         in_data[610],
                         in_data[729],
                         in_data[404],
                         in_data[581],
                         in_data[21],
                         in_data[203]
                    }),
            .out_data(lut_221_out)
        );

reg   lut_221_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_221_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_221_ff <= lut_221_out;
    end
end

assign out_data[221] = lut_221_ff;




// LUT : 222

wire lut_222_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001000110010111001101011100001101000100001001111001010111010),
            .DEVICE(DEVICE)
        )
    i_lut_222
        (
            .in_data({
                         in_data[2],
                         in_data[782],
                         in_data[537],
                         in_data[374],
                         in_data[772],
                         in_data[17]
                    }),
            .out_data(lut_222_out)
        );

reg   lut_222_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_222_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_222_ff <= lut_222_out;
    end
end

assign out_data[222] = lut_222_ff;




// LUT : 223

wire lut_223_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111111111010011110001111101011100011111110100110011111111010),
            .DEVICE(DEVICE)
        )
    i_lut_223
        (
            .in_data({
                         in_data[663],
                         in_data[397],
                         in_data[701],
                         in_data[425],
                         in_data[368],
                         in_data[430]
                    }),
            .out_data(lut_223_out)
        );

reg   lut_223_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_223_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_223_ff <= lut_223_out;
    end
end

assign out_data[223] = lut_223_ff;




// LUT : 224

wire lut_224_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111111111111011010110000111011111111001100110010101100001000),
            .DEVICE(DEVICE)
        )
    i_lut_224
        (
            .in_data({
                         in_data[270],
                         in_data[746],
                         in_data[495],
                         in_data[661],
                         in_data[699],
                         in_data[411]
                    }),
            .out_data(lut_224_out)
        );

reg   lut_224_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_224_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_224_ff <= lut_224_out;
    end
end

assign out_data[224] = lut_224_ff;




// LUT : 225

wire lut_225_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001001111010111110110011111100001111010111111101010011011001110),
            .DEVICE(DEVICE)
        )
    i_lut_225
        (
            .in_data({
                         in_data[715],
                         in_data[633],
                         in_data[609],
                         in_data[389],
                         in_data[733],
                         in_data[657]
                    }),
            .out_data(lut_225_out)
        );

reg   lut_225_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_225_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_225_ff <= lut_225_out;
    end
end

assign out_data[225] = lut_225_ff;




// LUT : 226

wire lut_226_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101001001110101000001000001011101110110010101010101011010000),
            .DEVICE(DEVICE)
        )
    i_lut_226
        (
            .in_data({
                         in_data[492],
                         in_data[69],
                         in_data[601],
                         in_data[571],
                         in_data[189],
                         in_data[731]
                    }),
            .out_data(lut_226_out)
        );

reg   lut_226_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_226_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_226_ff <= lut_226_out;
    end
end

assign out_data[226] = lut_226_ff;




// LUT : 227

wire lut_227_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101001010100110110110101101011101010010111100101011111011110100),
            .DEVICE(DEVICE)
        )
    i_lut_227
        (
            .in_data({
                         in_data[248],
                         in_data[472],
                         in_data[470],
                         in_data[777],
                         in_data[616],
                         in_data[704]
                    }),
            .out_data(lut_227_out)
        );

reg   lut_227_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_227_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_227_ff <= lut_227_out;
    end
end

assign out_data[227] = lut_227_ff;




// LUT : 228

wire lut_228_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111001001111101000010101001000111100110001001010000011110010111),
            .DEVICE(DEVICE)
        )
    i_lut_228
        (
            .in_data({
                         in_data[522],
                         in_data[447],
                         in_data[217],
                         in_data[286],
                         in_data[185],
                         in_data[737]
                    }),
            .out_data(lut_228_out)
        );

reg   lut_228_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_228_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_228_ff <= lut_228_out;
    end
end

assign out_data[228] = lut_228_ff;




// LUT : 229

wire lut_229_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111001110001010000011001111010101101000000000110010100111010),
            .DEVICE(DEVICE)
        )
    i_lut_229
        (
            .in_data({
                         in_data[734],
                         in_data[345],
                         in_data[5],
                         in_data[242],
                         in_data[665],
                         in_data[666]
                    }),
            .out_data(lut_229_out)
        );

reg   lut_229_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_229_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_229_ff <= lut_229_out;
    end
end

assign out_data[229] = lut_229_ff;




// LUT : 230

wire lut_230_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101011010110010110111001001110101000001111100111101110000000),
            .DEVICE(DEVICE)
        )
    i_lut_230
        (
            .in_data({
                         in_data[543],
                         in_data[6],
                         in_data[156],
                         in_data[298],
                         in_data[56],
                         in_data[177]
                    }),
            .out_data(lut_230_out)
        );

reg   lut_230_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_230_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_230_ff <= lut_230_out;
    end
end

assign out_data[230] = lut_230_ff;




// LUT : 231

wire lut_231_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011010111100110000011111001111110110010011001011111101001100),
            .DEVICE(DEVICE)
        )
    i_lut_231
        (
            .in_data({
                         in_data[250],
                         in_data[310],
                         in_data[99],
                         in_data[681],
                         in_data[559],
                         in_data[157]
                    }),
            .out_data(lut_231_out)
        );

reg   lut_231_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_231_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_231_ff <= lut_231_out;
    end
end

assign out_data[231] = lut_231_ff;




// LUT : 232

wire lut_232_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000111011011110010100101101000110110100001101010000111011111),
            .DEVICE(DEVICE)
        )
    i_lut_232
        (
            .in_data({
                         in_data[381],
                         in_data[392],
                         in_data[361],
                         in_data[34],
                         in_data[654],
                         in_data[675]
                    }),
            .out_data(lut_232_out)
        );

reg   lut_232_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_232_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_232_ff <= lut_232_out;
    end
end

assign out_data[232] = lut_232_ff;




// LUT : 233

wire lut_233_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110110001010010100100101010101110001000010000001101011101000000),
            .DEVICE(DEVICE)
        )
    i_lut_233
        (
            .in_data({
                         in_data[450],
                         in_data[62],
                         in_data[296],
                         in_data[258],
                         in_data[369],
                         in_data[370]
                    }),
            .out_data(lut_233_out)
        );

reg   lut_233_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_233_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_233_ff <= lut_233_out;
    end
end

assign out_data[233] = lut_233_ff;




// LUT : 234

wire lut_234_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001001000100010001000001011001110101010101011011010100110101),
            .DEVICE(DEVICE)
        )
    i_lut_234
        (
            .in_data({
                         in_data[639],
                         in_data[128],
                         in_data[271],
                         in_data[783],
                         in_data[732],
                         in_data[251]
                    }),
            .out_data(lut_234_out)
        );

reg   lut_234_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_234_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_234_ff <= lut_234_out;
    end
end

assign out_data[234] = lut_234_ff;




// LUT : 235

wire lut_235_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101001110000101111111011111110111010111100111111111111111111101),
            .DEVICE(DEVICE)
        )
    i_lut_235
        (
            .in_data({
                         in_data[490],
                         in_data[92],
                         in_data[293],
                         in_data[719],
                         in_data[232],
                         in_data[351]
                    }),
            .out_data(lut_235_out)
        );

reg   lut_235_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_235_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_235_ff <= lut_235_out;
    end
end

assign out_data[235] = lut_235_ff;




// LUT : 236

wire lut_236_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001100111001111100011011100110010010001011101010010011100100),
            .DEVICE(DEVICE)
        )
    i_lut_236
        (
            .in_data({
                         in_data[47],
                         in_data[426],
                         in_data[362],
                         in_data[132],
                         in_data[658],
                         in_data[284]
                    }),
            .out_data(lut_236_out)
        );

reg   lut_236_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_236_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_236_ff <= lut_236_out;
    end
end

assign out_data[236] = lut_236_ff;




// LUT : 237

wire lut_237_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010110001000011001000000100010010001110011011110100000011001),
            .DEVICE(DEVICE)
        )
    i_lut_237
        (
            .in_data({
                         in_data[508],
                         in_data[181],
                         in_data[645],
                         in_data[595],
                         in_data[403],
                         in_data[429]
                    }),
            .out_data(lut_237_out)
        );

reg   lut_237_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_237_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_237_ff <= lut_237_out;
    end
end

assign out_data[237] = lut_237_ff;




// LUT : 238

wire lut_238_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001000111010111101001101011000100011100000101111110001111101),
            .DEVICE(DEVICE)
        )
    i_lut_238
        (
            .in_data({
                         in_data[680],
                         in_data[423],
                         in_data[740],
                         in_data[596],
                         in_data[622],
                         in_data[33]
                    }),
            .out_data(lut_238_out)
        );

reg   lut_238_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_238_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_238_ff <= lut_238_out;
    end
end

assign out_data[238] = lut_238_ff;




// LUT : 239

wire lut_239_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100010111001011110001000111001000111011010011000110111000100010),
            .DEVICE(DEVICE)
        )
    i_lut_239
        (
            .in_data({
                         in_data[691],
                         in_data[14],
                         in_data[676],
                         in_data[231],
                         in_data[424],
                         in_data[249]
                    }),
            .out_data(lut_239_out)
        );

reg   lut_239_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_239_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_239_ff <= lut_239_out;
    end
end

assign out_data[239] = lut_239_ff;




// LUT : 240

wire lut_240_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101100100111000001010000010110011111001110000000010000000100),
            .DEVICE(DEVICE)
        )
    i_lut_240
        (
            .in_data({
                         in_data[526],
                         in_data[685],
                         in_data[579],
                         in_data[377],
                         in_data[499],
                         in_data[96]
                    }),
            .out_data(lut_240_out)
        );

reg   lut_240_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_240_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_240_ff <= lut_240_out;
    end
end

assign out_data[240] = lut_240_ff;




// LUT : 241

wire lut_241_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111101000000000000000110110000110001000000100110000010000010),
            .DEVICE(DEVICE)
        )
    i_lut_241
        (
            .in_data({
                         in_data[130],
                         in_data[435],
                         in_data[512],
                         in_data[238],
                         in_data[61],
                         in_data[532]
                    }),
            .out_data(lut_241_out)
        );

reg   lut_241_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_241_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_241_ff <= lut_241_out;
    end
end

assign out_data[241] = lut_241_ff;




// LUT : 242

wire lut_242_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000010011100100010101110100010010110001001000001110000000000),
            .DEVICE(DEVICE)
        )
    i_lut_242
        (
            .in_data({
                         in_data[182],
                         in_data[198],
                         in_data[629],
                         in_data[41],
                         in_data[48],
                         in_data[754]
                    }),
            .out_data(lut_242_out)
        );

reg   lut_242_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_242_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_242_ff <= lut_242_out;
    end
end

assign out_data[242] = lut_242_ff;




// LUT : 243

wire lut_243_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110100011110100001010110111111011001110001110001000011011111),
            .DEVICE(DEVICE)
        )
    i_lut_243
        (
            .in_data({
                         in_data[556],
                         in_data[282],
                         in_data[54],
                         in_data[109],
                         in_data[211],
                         in_data[529]
                    }),
            .out_data(lut_243_out)
        );

reg   lut_243_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_243_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_243_ff <= lut_243_out;
    end
end

assign out_data[243] = lut_243_ff;




// LUT : 244

wire lut_244_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110011101111010111001111111101111111100011001100111101001100),
            .DEVICE(DEVICE)
        )
    i_lut_244
        (
            .in_data({
                         in_data[528],
                         in_data[215],
                         in_data[591],
                         in_data[288],
                         in_data[611],
                         in_data[630]
                    }),
            .out_data(lut_244_out)
        );

reg   lut_244_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_244_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_244_ff <= lut_244_out;
    end
end

assign out_data[244] = lut_244_ff;




// LUT : 245

wire lut_245_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111011111011110010101000100110000010100000101000100110000101),
            .DEVICE(DEVICE)
        )
    i_lut_245
        (
            .in_data({
                         in_data[317],
                         in_data[781],
                         in_data[83],
                         in_data[723],
                         in_data[563],
                         in_data[692]
                    }),
            .out_data(lut_245_out)
        );

reg   lut_245_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_245_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_245_ff <= lut_245_out;
    end
end

assign out_data[245] = lut_245_ff;




// LUT : 246

wire lut_246_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111110101111000100110111111100110001101001011000001101110001),
            .DEVICE(DEVICE)
        )
    i_lut_246
        (
            .in_data({
                         in_data[409],
                         in_data[688],
                         in_data[684],
                         in_data[334],
                         in_data[87],
                         in_data[243]
                    }),
            .out_data(lut_246_out)
        );

reg   lut_246_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_246_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_246_ff <= lut_246_out;
    end
end

assign out_data[246] = lut_246_ff;




// LUT : 247

wire lut_247_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110010010010101101011100111001100111111001111001111011001110),
            .DEVICE(DEVICE)
        )
    i_lut_247
        (
            .in_data({
                         in_data[247],
                         in_data[474],
                         in_data[642],
                         in_data[340],
                         in_data[212],
                         in_data[780]
                    }),
            .out_data(lut_247_out)
        );

reg   lut_247_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_247_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_247_ff <= lut_247_out;
    end
end

assign out_data[247] = lut_247_ff;




// LUT : 248

wire lut_248_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010101011011011101011111011100010111011011111001011100101001),
            .DEVICE(DEVICE)
        )
    i_lut_248
        (
            .in_data({
                         in_data[523],
                         in_data[318],
                         in_data[311],
                         in_data[338],
                         in_data[86],
                         in_data[91]
                    }),
            .out_data(lut_248_out)
        );

reg   lut_248_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_248_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_248_ff <= lut_248_out;
    end
end

assign out_data[248] = lut_248_ff;




// LUT : 249

wire lut_249_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101001111010011110001010100000001100001000001111101100010001),
            .DEVICE(DEVICE)
        )
    i_lut_249
        (
            .in_data({
                         in_data[225],
                         in_data[418],
                         in_data[720],
                         in_data[358],
                         in_data[279],
                         in_data[72]
                    }),
            .out_data(lut_249_out)
        );

reg   lut_249_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_249_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_249_ff <= lut_249_out;
    end
end

assign out_data[249] = lut_249_ff;




// LUT : 250

wire lut_250_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000010111111110101111110011110100101011010011101111100101010),
            .DEVICE(DEVICE)
        )
    i_lut_250
        (
            .in_data({
                         in_data[627],
                         in_data[502],
                         in_data[749],
                         in_data[60],
                         in_data[356],
                         in_data[256]
                    }),
            .out_data(lut_250_out)
        );

reg   lut_250_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_250_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_250_ff <= lut_250_out;
    end
end

assign out_data[250] = lut_250_ff;




// LUT : 251

wire lut_251_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110011110101101100110111010110011111010111000101000101010100),
            .DEVICE(DEVICE)
        )
    i_lut_251
        (
            .in_data({
                         in_data[202],
                         in_data[384],
                         in_data[11],
                         in_data[469],
                         in_data[586],
                         in_data[770]
                    }),
            .out_data(lut_251_out)
        );

reg   lut_251_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_251_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_251_ff <= lut_251_out;
    end
end

assign out_data[251] = lut_251_ff;




// LUT : 252

wire lut_252_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010110111100011111101010010100111111110011110010001001010111),
            .DEVICE(DEVICE)
        )
    i_lut_252
        (
            .in_data({
                         in_data[448],
                         in_data[37],
                         in_data[287],
                         in_data[631],
                         in_data[199],
                         in_data[280]
                    }),
            .out_data(lut_252_out)
        );

reg   lut_252_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_252_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_252_ff <= lut_252_out;
    end
end

assign out_data[252] = lut_252_ff;




// LUT : 253

wire lut_253_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000111001010110110101100111110100101010101011111111011000000),
            .DEVICE(DEVICE)
        )
    i_lut_253
        (
            .in_data({
                         in_data[200],
                         in_data[728],
                         in_data[518],
                         in_data[193],
                         in_data[333],
                         in_data[292]
                    }),
            .out_data(lut_253_out)
        );

reg   lut_253_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_253_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_253_ff <= lut_253_out;
    end
end

assign out_data[253] = lut_253_ff;




// LUT : 254

wire lut_254_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101111001000100011010110000010000111110010001101000100110000),
            .DEVICE(DEVICE)
        )
    i_lut_254
        (
            .in_data({
                         in_data[295],
                         in_data[108],
                         in_data[709],
                         in_data[565],
                         in_data[752],
                         in_data[541]
                    }),
            .out_data(lut_254_out)
        );

reg   lut_254_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_254_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_254_ff <= lut_254_out;
    end
end

assign out_data[254] = lut_254_ff;




// LUT : 255

wire lut_255_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000100010010101000011111011110101010010111111110101000010101),
            .DEVICE(DEVICE)
        )
    i_lut_255
        (
            .in_data({
                         in_data[449],
                         in_data[483],
                         in_data[441],
                         in_data[511],
                         in_data[184],
                         in_data[664]
                    }),
            .out_data(lut_255_out)
        );

reg   lut_255_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_255_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_255_ff <= lut_255_out;
    end
end

assign out_data[255] = lut_255_ff;




// LUT : 256

wire lut_256_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001110100101000100110000000010101100110110000100001101011011),
            .DEVICE(DEVICE)
        )
    i_lut_256
        (
            .in_data({
                         in_data[4],
                         in_data[104],
                         in_data[707],
                         in_data[530],
                         in_data[102],
                         in_data[761]
                    }),
            .out_data(lut_256_out)
        );

reg   lut_256_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_256_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_256_ff <= lut_256_out;
    end
end

assign out_data[256] = lut_256_ff;




// LUT : 257

wire lut_257_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110111111111110011001110101011101000101001000100000000001100),
            .DEVICE(DEVICE)
        )
    i_lut_257
        (
            .in_data({
                         in_data[71],
                         in_data[741],
                         in_data[233],
                         in_data[582],
                         in_data[28],
                         in_data[456]
                    }),
            .out_data(lut_257_out)
        );

reg   lut_257_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_257_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_257_ff <= lut_257_out;
    end
end

assign out_data[257] = lut_257_ff;




// LUT : 258

wire lut_258_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101100001111010110001111101011001001000110000001010000000101110),
            .DEVICE(DEVICE)
        )
    i_lut_258
        (
            .in_data({
                         in_data[140],
                         in_data[673],
                         in_data[558],
                         in_data[39],
                         in_data[214],
                         in_data[31]
                    }),
            .out_data(lut_258_out)
        );

reg   lut_258_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_258_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_258_ff <= lut_258_out;
    end
end

assign out_data[258] = lut_258_ff;




// LUT : 259

wire lut_259_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111110001111011101100011011111100110100010100011010011110110),
            .DEVICE(DEVICE)
        )
    i_lut_259
        (
            .in_data({
                         in_data[235],
                         in_data[164],
                         in_data[710],
                         in_data[278],
                         in_data[717],
                         in_data[548]
                    }),
            .out_data(lut_259_out)
        );

reg   lut_259_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_259_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_259_ff <= lut_259_out;
    end
end

assign out_data[259] = lut_259_ff;




// LUT : 260

wire lut_260_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101010110000101001110110111101100101011001111111110101111001),
            .DEVICE(DEVICE)
        )
    i_lut_260
        (
            .in_data({
                         in_data[43],
                         in_data[103],
                         in_data[487],
                         in_data[705],
                         in_data[569],
                         in_data[168]
                    }),
            .out_data(lut_260_out)
        );

reg   lut_260_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_260_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_260_ff <= lut_260_out;
    end
end

assign out_data[260] = lut_260_ff;




// LUT : 261

wire lut_261_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011101000010000010000000010101000100111110100000001011000100),
            .DEVICE(DEVICE)
        )
    i_lut_261
        (
            .in_data({
                         in_data[295],
                         in_data[668],
                         in_data[220],
                         in_data[529],
                         in_data[267],
                         in_data[70]
                    }),
            .out_data(lut_261_out)
        );

reg   lut_261_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_261_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_261_ff <= lut_261_out;
    end
end

assign out_data[261] = lut_261_ff;




// LUT : 262

wire lut_262_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100010111110011101111100111010011111101110001000101010100000000),
            .DEVICE(DEVICE)
        )
    i_lut_262
        (
            .in_data({
                         in_data[16],
                         in_data[161],
                         in_data[235],
                         in_data[602],
                         in_data[303],
                         in_data[541]
                    }),
            .out_data(lut_262_out)
        );

reg   lut_262_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_262_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_262_ff <= lut_262_out;
    end
end

assign out_data[262] = lut_262_ff;




// LUT : 263

wire lut_263_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010100001111111011110010011100011100010101010100000100001001),
            .DEVICE(DEVICE)
        )
    i_lut_263
        (
            .in_data({
                         in_data[479],
                         in_data[87],
                         in_data[150],
                         in_data[727],
                         in_data[408],
                         in_data[737]
                    }),
            .out_data(lut_263_out)
        );

reg   lut_263_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_263_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_263_ff <= lut_263_out;
    end
end

assign out_data[263] = lut_263_ff;




// LUT : 264

wire lut_264_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010100111111010111011111011110100111110011111001111101111000),
            .DEVICE(DEVICE)
        )
    i_lut_264
        (
            .in_data({
                         in_data[297],
                         in_data[642],
                         in_data[556],
                         in_data[459],
                         in_data[441],
                         in_data[421]
                    }),
            .out_data(lut_264_out)
        );

reg   lut_264_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_264_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_264_ff <= lut_264_out;
    end
end

assign out_data[264] = lut_264_ff;




// LUT : 265

wire lut_265_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111111010101111100010000111001101001000010000101010100110001),
            .DEVICE(DEVICE)
        )
    i_lut_265
        (
            .in_data({
                         in_data[694],
                         in_data[107],
                         in_data[473],
                         in_data[600],
                         in_data[733],
                         in_data[57]
                    }),
            .out_data(lut_265_out)
        );

reg   lut_265_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_265_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_265_ff <= lut_265_out;
    end
end

assign out_data[265] = lut_265_ff;




// LUT : 266

wire lut_266_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101000101110000001111000000000010011100000001011011100101011),
            .DEVICE(DEVICE)
        )
    i_lut_266
        (
            .in_data({
                         in_data[690],
                         in_data[632],
                         in_data[587],
                         in_data[423],
                         in_data[469],
                         in_data[588]
                    }),
            .out_data(lut_266_out)
        );

reg   lut_266_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_266_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_266_ff <= lut_266_out;
    end
end

assign out_data[266] = lut_266_ff;




// LUT : 267

wire lut_267_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110001101000101011001011100001000100110011001000011111001101),
            .DEVICE(DEVICE)
        )
    i_lut_267
        (
            .in_data({
                         in_data[164],
                         in_data[597],
                         in_data[346],
                         in_data[79],
                         in_data[59],
                         in_data[240]
                    }),
            .out_data(lut_267_out)
        );

reg   lut_267_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_267_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_267_ff <= lut_267_out;
    end
end

assign out_data[267] = lut_267_ff;




// LUT : 268

wire lut_268_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000110111100101100111000000101011001001000100011101100000100),
            .DEVICE(DEVICE)
        )
    i_lut_268
        (
            .in_data({
                         in_data[717],
                         in_data[503],
                         in_data[641],
                         in_data[686],
                         in_data[679],
                         in_data[306]
                    }),
            .out_data(lut_268_out)
        );

reg   lut_268_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_268_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_268_ff <= lut_268_out;
    end
end

assign out_data[268] = lut_268_ff;




// LUT : 269

wire lut_269_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001101111111001101001110110001111010011101111011111111111100),
            .DEVICE(DEVICE)
        )
    i_lut_269
        (
            .in_data({
                         in_data[552],
                         in_data[144],
                         in_data[222],
                         in_data[596],
                         in_data[121],
                         in_data[291]
                    }),
            .out_data(lut_269_out)
        );

reg   lut_269_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_269_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_269_ff <= lut_269_out;
    end
end

assign out_data[269] = lut_269_ff;




// LUT : 270

wire lut_270_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001101000000000100110100001110100101000111010101100100000100000),
            .DEVICE(DEVICE)
        )
    i_lut_270
        (
            .in_data({
                         in_data[286],
                         in_data[230],
                         in_data[464],
                         in_data[615],
                         in_data[661],
                         in_data[8]
                    }),
            .out_data(lut_270_out)
        );

reg   lut_270_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_270_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_270_ff <= lut_270_out;
    end
end

assign out_data[270] = lut_270_ff;




// LUT : 271

wire lut_271_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110000101011000100010110001110001011010110101110110001000100),
            .DEVICE(DEVICE)
        )
    i_lut_271
        (
            .in_data({
                         in_data[532],
                         in_data[45],
                         in_data[47],
                         in_data[652],
                         in_data[765],
                         in_data[125]
                    }),
            .out_data(lut_271_out)
        );

reg   lut_271_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_271_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_271_ff <= lut_271_out;
    end
end

assign out_data[271] = lut_271_ff;




// LUT : 272

wire lut_272_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000011110001110100100000101000000000101000111111),
            .DEVICE(DEVICE)
        )
    i_lut_272
        (
            .in_data({
                         in_data[659],
                         in_data[380],
                         in_data[126],
                         in_data[320],
                         in_data[205],
                         in_data[315]
                    }),
            .out_data(lut_272_out)
        );

reg   lut_272_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_272_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_272_ff <= lut_272_out;
    end
end

assign out_data[272] = lut_272_ff;




// LUT : 273

wire lut_273_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011110011110111111000011111011111000110111111000101011011101110),
            .DEVICE(DEVICE)
        )
    i_lut_273
        (
            .in_data({
                         in_data[611],
                         in_data[257],
                         in_data[756],
                         in_data[187],
                         in_data[623],
                         in_data[284]
                    }),
            .out_data(lut_273_out)
        );

reg   lut_273_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_273_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_273_ff <= lut_273_out;
    end
end

assign out_data[273] = lut_273_ff;




// LUT : 274

wire lut_274_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010100010101100101011101000111011010011001101111100101110000),
            .DEVICE(DEVICE)
        )
    i_lut_274
        (
            .in_data({
                         in_data[329],
                         in_data[171],
                         in_data[64],
                         in_data[343],
                         in_data[130],
                         in_data[365]
                    }),
            .out_data(lut_274_out)
        );

reg   lut_274_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_274_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_274_ff <= lut_274_out;
    end
end

assign out_data[274] = lut_274_ff;




// LUT : 275

wire lut_275_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001010001101010110001110111011100001011101110111010001110011),
            .DEVICE(DEVICE)
        )
    i_lut_275
        (
            .in_data({
                         in_data[111],
                         in_data[713],
                         in_data[35],
                         in_data[631],
                         in_data[75],
                         in_data[154]
                    }),
            .out_data(lut_275_out)
        );

reg   lut_275_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_275_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_275_ff <= lut_275_out;
    end
end

assign out_data[275] = lut_275_ff;




// LUT : 276

wire lut_276_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101100000111010000111010100010111111011000000110001100010101010),
            .DEVICE(DEVICE)
        )
    i_lut_276
        (
            .in_data({
                         in_data[224],
                         in_data[772],
                         in_data[78],
                         in_data[557],
                         in_data[751],
                         in_data[714]
                    }),
            .out_data(lut_276_out)
        );

reg   lut_276_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_276_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_276_ff <= lut_276_out;
    end
end

assign out_data[276] = lut_276_ff;




// LUT : 277

wire lut_277_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110011101000101010101001000010010010111101011101001011110111),
            .DEVICE(DEVICE)
        )
    i_lut_277
        (
            .in_data({
                         in_data[173],
                         in_data[292],
                         in_data[116],
                         in_data[501],
                         in_data[715],
                         in_data[31]
                    }),
            .out_data(lut_277_out)
        );

reg   lut_277_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_277_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_277_ff <= lut_277_out;
    end
end

assign out_data[277] = lut_277_ff;




// LUT : 278

wire lut_278_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010101010001110000111110110010101000101000011010001111010001),
            .DEVICE(DEVICE)
        )
    i_lut_278
        (
            .in_data({
                         in_data[310],
                         in_data[766],
                         in_data[102],
                         in_data[530],
                         in_data[534],
                         in_data[630]
                    }),
            .out_data(lut_278_out)
        );

reg   lut_278_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_278_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_278_ff <= lut_278_out;
    end
end

assign out_data[278] = lut_278_ff;




// LUT : 279

wire lut_279_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001101011110101000010001111000011110010010111001111111011111110),
            .DEVICE(DEVICE)
        )
    i_lut_279
        (
            .in_data({
                         in_data[85],
                         in_data[709],
                         in_data[438],
                         in_data[434],
                         in_data[542],
                         in_data[95]
                    }),
            .out_data(lut_279_out)
        );

reg   lut_279_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_279_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_279_ff <= lut_279_out;
    end
end

assign out_data[279] = lut_279_ff;




// LUT : 280

wire lut_280_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010010110010010011111110111001100110101010101010011111101111),
            .DEVICE(DEVICE)
        )
    i_lut_280
        (
            .in_data({
                         in_data[182],
                         in_data[720],
                         in_data[90],
                         in_data[159],
                         in_data[323],
                         in_data[340]
                    }),
            .out_data(lut_280_out)
        );

reg   lut_280_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_280_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_280_ff <= lut_280_out;
    end
end

assign out_data[280] = lut_280_ff;




// LUT : 281

wire lut_281_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111100101110001000001010010010101111000011001010001000001101),
            .DEVICE(DEVICE)
        )
    i_lut_281
        (
            .in_data({
                         in_data[158],
                         in_data[215],
                         in_data[129],
                         in_data[276],
                         in_data[513],
                         in_data[314]
                    }),
            .out_data(lut_281_out)
        );

reg   lut_281_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_281_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_281_ff <= lut_281_out;
    end
end

assign out_data[281] = lut_281_ff;




// LUT : 282

wire lut_282_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101100001011000110110110111111000000010110010000000001111000),
            .DEVICE(DEVICE)
        )
    i_lut_282
        (
            .in_data({
                         in_data[305],
                         in_data[410],
                         in_data[127],
                         in_data[767],
                         in_data[551],
                         in_data[476]
                    }),
            .out_data(lut_282_out)
        );

reg   lut_282_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_282_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_282_ff <= lut_282_out;
    end
end

assign out_data[282] = lut_282_ff;




// LUT : 283

wire lut_283_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100110000110011011010001000101000100000001000011000011010101),
            .DEVICE(DEVICE)
        )
    i_lut_283
        (
            .in_data({
                         in_data[65],
                         in_data[321],
                         in_data[625],
                         in_data[175],
                         in_data[312],
                         in_data[570]
                    }),
            .out_data(lut_283_out)
        );

reg   lut_283_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_283_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_283_ff <= lut_283_out;
    end
end

assign out_data[283] = lut_283_ff;




// LUT : 284

wire lut_284_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111110011111001100110100000011001000111011101111010001100101111),
            .DEVICE(DEVICE)
        )
    i_lut_284
        (
            .in_data({
                         in_data[356],
                         in_data[392],
                         in_data[658],
                         in_data[695],
                         in_data[169],
                         in_data[418]
                    }),
            .out_data(lut_284_out)
        );

reg   lut_284_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_284_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_284_ff <= lut_284_out;
    end
end

assign out_data[284] = lut_284_ff;




// LUT : 285

wire lut_285_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101110001010110011001010000011001100110111110110001100100011),
            .DEVICE(DEVICE)
        )
    i_lut_285
        (
            .in_data({
                         in_data[782],
                         in_data[443],
                         in_data[375],
                         in_data[477],
                         in_data[378],
                         in_data[298]
                    }),
            .out_data(lut_285_out)
        );

reg   lut_285_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_285_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_285_ff <= lut_285_out;
    end
end

assign out_data[285] = lut_285_ff;




// LUT : 286

wire lut_286_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000110010001011001000111110111100011111101011011100100110000),
            .DEVICE(DEVICE)
        )
    i_lut_286
        (
            .in_data({
                         in_data[219],
                         in_data[653],
                         in_data[81],
                         in_data[462],
                         in_data[497],
                         in_data[417]
                    }),
            .out_data(lut_286_out)
        );

reg   lut_286_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_286_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_286_ff <= lut_286_out;
    end
end

assign out_data[286] = lut_286_ff;




// LUT : 287

wire lut_287_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001101101110111100110111111010111001001001100111011111110110),
            .DEVICE(DEVICE)
        )
    i_lut_287
        (
            .in_data({
                         in_data[680],
                         in_data[638],
                         in_data[424],
                         in_data[377],
                         in_data[254],
                         in_data[708]
                    }),
            .out_data(lut_287_out)
        );

reg   lut_287_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_287_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_287_ff <= lut_287_out;
    end
end

assign out_data[287] = lut_287_ff;




// LUT : 288

wire lut_288_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001101000100100001010000000001011010111100011001000110000101010),
            .DEVICE(DEVICE)
        )
    i_lut_288
        (
            .in_data({
                         in_data[707],
                         in_data[283],
                         in_data[616],
                         in_data[579],
                         in_data[669],
                         in_data[316]
                    }),
            .out_data(lut_288_out)
        );

reg   lut_288_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_288_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_288_ff <= lut_288_out;
    end
end

assign out_data[288] = lut_288_ff;




// LUT : 289

wire lut_289_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011011100110001010000001100011100101001000010100100101001011),
            .DEVICE(DEVICE)
        )
    i_lut_289
        (
            .in_data({
                         in_data[190],
                         in_data[736],
                         in_data[133],
                         in_data[366],
                         in_data[391],
                         in_data[98]
                    }),
            .out_data(lut_289_out)
        );

reg   lut_289_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_289_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_289_ff <= lut_289_out;
    end
end

assign out_data[289] = lut_289_ff;




// LUT : 290

wire lut_290_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111100101111010111101110101010111111100010101110101011011010),
            .DEVICE(DEVICE)
        )
    i_lut_290
        (
            .in_data({
                         in_data[660],
                         in_data[155],
                         in_data[406],
                         in_data[3],
                         in_data[275],
                         in_data[201]
                    }),
            .out_data(lut_290_out)
        );

reg   lut_290_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_290_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_290_ff <= lut_290_out;
    end
end

assign out_data[290] = lut_290_ff;




// LUT : 291

wire lut_291_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100001010010011011110000011110110010100000100100111001000111),
            .DEVICE(DEVICE)
        )
    i_lut_291
        (
            .in_data({
                         in_data[577],
                         in_data[143],
                         in_data[496],
                         in_data[99],
                         in_data[231],
                         in_data[132]
                    }),
            .out_data(lut_291_out)
        );

reg   lut_291_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_291_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_291_ff <= lut_291_out;
    end
end

assign out_data[291] = lut_291_ff;




// LUT : 292

wire lut_292_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001110001010001110001001000011001000101100000111001111000001),
            .DEVICE(DEVICE)
        )
    i_lut_292
        (
            .in_data({
                         in_data[247],
                         in_data[337],
                         in_data[165],
                         in_data[141],
                         in_data[735],
                         in_data[711]
                    }),
            .out_data(lut_292_out)
        );

reg   lut_292_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_292_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_292_ff <= lut_292_out;
    end
end

assign out_data[292] = lut_292_ff;




// LUT : 293

wire lut_293_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000100001111101111001101100001011000111101011011110011110111110),
            .DEVICE(DEVICE)
        )
    i_lut_293
        (
            .in_data({
                         in_data[516],
                         in_data[71],
                         in_data[53],
                         in_data[505],
                         in_data[307],
                         in_data[774]
                    }),
            .out_data(lut_293_out)
        );

reg   lut_293_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_293_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_293_ff <= lut_293_out;
    end
end

assign out_data[293] = lut_293_ff;




// LUT : 294

wire lut_294_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010011101101000010000000100100011110011011111111111010010000100),
            .DEVICE(DEVICE)
        )
    i_lut_294
        (
            .in_data({
                         in_data[397],
                         in_data[543],
                         in_data[522],
                         in_data[635],
                         in_data[672],
                         in_data[273]
                    }),
            .out_data(lut_294_out)
        );

reg   lut_294_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_294_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_294_ff <= lut_294_out;
    end
end

assign out_data[294] = lut_294_ff;




// LUT : 295

wire lut_295_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001101101001011110000000110100000101000110010100100001001),
            .DEVICE(DEVICE)
        )
    i_lut_295
        (
            .in_data({
                         in_data[467],
                         in_data[637],
                         in_data[608],
                         in_data[260],
                         in_data[194],
                         in_data[704]
                    }),
            .out_data(lut_295_out)
        );

reg   lut_295_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_295_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_295_ff <= lut_295_out;
    end
end

assign out_data[295] = lut_295_ff;




// LUT : 296

wire lut_296_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010111001101101110010100011100010101011010011000000101010001110),
            .DEVICE(DEVICE)
        )
    i_lut_296
        (
            .in_data({
                         in_data[644],
                         in_data[341],
                         in_data[678],
                         in_data[289],
                         in_data[269],
                         in_data[429]
                    }),
            .out_data(lut_296_out)
        );

reg   lut_296_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_296_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_296_ff <= lut_296_out;
    end
end

assign out_data[296] = lut_296_ff;




// LUT : 297

wire lut_297_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111110010110011010000010101000110110111100101100010011110000),
            .DEVICE(DEVICE)
        )
    i_lut_297
        (
            .in_data({
                         in_data[309],
                         in_data[91],
                         in_data[367],
                         in_data[350],
                         in_data[547],
                         in_data[629]
                    }),
            .out_data(lut_297_out)
        );

reg   lut_297_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_297_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_297_ff <= lut_297_out;
    end
end

assign out_data[297] = lut_297_ff;




// LUT : 298

wire lut_298_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110011010011101000001011011110111110100111111001011101110101010),
            .DEVICE(DEVICE)
        )
    i_lut_298
        (
            .in_data({
                         in_data[393],
                         in_data[56],
                         in_data[622],
                         in_data[436],
                         in_data[294],
                         in_data[639]
                    }),
            .out_data(lut_298_out)
        );

reg   lut_298_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_298_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_298_ff <= lut_298_out;
    end
end

assign out_data[298] = lut_298_ff;




// LUT : 299

wire lut_299_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110000001011110010001011011011101101111101111010110011110101),
            .DEVICE(DEVICE)
        )
    i_lut_299
        (
            .in_data({
                         in_data[673],
                         in_data[262],
                         in_data[728],
                         in_data[279],
                         in_data[521],
                         in_data[352]
                    }),
            .out_data(lut_299_out)
        );

reg   lut_299_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_299_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_299_ff <= lut_299_out;
    end
end

assign out_data[299] = lut_299_ff;




// LUT : 300

wire lut_300_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111001111101011100010000101101100001110011011000101111101011),
            .DEVICE(DEVICE)
        )
    i_lut_300
        (
            .in_data({
                         in_data[131],
                         in_data[399],
                         in_data[757],
                         in_data[665],
                         in_data[583],
                         in_data[750]
                    }),
            .out_data(lut_300_out)
        );

reg   lut_300_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_300_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_300_ff <= lut_300_out;
    end
end

assign out_data[300] = lut_300_ff;




// LUT : 301

wire lut_301_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110001111111001101111111001010000010100010100111010101111011),
            .DEVICE(DEVICE)
        )
    i_lut_301
        (
            .in_data({
                         in_data[390],
                         in_data[22],
                         in_data[243],
                         in_data[191],
                         in_data[490],
                         in_data[72]
                    }),
            .out_data(lut_301_out)
        );

reg   lut_301_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_301_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_301_ff <= lut_301_out;
    end
end

assign out_data[301] = lut_301_ff;




// LUT : 302

wire lut_302_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100000101011001011000100101001100111010100111011100100010001),
            .DEVICE(DEVICE)
        )
    i_lut_302
        (
            .in_data({
                         in_data[134],
                         in_data[396],
                         in_data[491],
                         in_data[318],
                         in_data[40],
                         in_data[363]
                    }),
            .out_data(lut_302_out)
        );

reg   lut_302_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_302_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_302_ff <= lut_302_out;
    end
end

assign out_data[302] = lut_302_ff;




// LUT : 303

wire lut_303_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101011001000000101000000000100100000101010100000111000101110),
            .DEVICE(DEVICE)
        )
    i_lut_303
        (
            .in_data({
                         in_data[761],
                         in_data[370],
                         in_data[688],
                         in_data[607],
                         in_data[234],
                         in_data[29]
                    }),
            .out_data(lut_303_out)
        );

reg   lut_303_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_303_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_303_ff <= lut_303_out;
    end
end

assign out_data[303] = lut_303_ff;




// LUT : 304

wire lut_304_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000011110000000000001110000001001100110100000000100111110101),
            .DEVICE(DEVICE)
        )
    i_lut_304
        (
            .in_data({
                         in_data[572],
                         in_data[302],
                         in_data[96],
                         in_data[416],
                         in_data[242],
                         in_data[357]
                    }),
            .out_data(lut_304_out)
        );

reg   lut_304_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_304_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_304_ff <= lut_304_out;
    end
end

assign out_data[304] = lut_304_ff;




// LUT : 305

wire lut_305_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010000111111000001101111111001110101001111111110110111110100),
            .DEVICE(DEVICE)
        )
    i_lut_305
        (
            .in_data({
                         in_data[682],
                         in_data[667],
                         in_data[189],
                         in_data[643],
                         in_data[666],
                         in_data[465]
                    }),
            .out_data(lut_305_out)
        );

reg   lut_305_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_305_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_305_ff <= lut_305_out;
    end
end

assign out_data[305] = lut_305_ff;




// LUT : 306

wire lut_306_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100000010111100001000011011100100000111110110111010010110011),
            .DEVICE(DEVICE)
        )
    i_lut_306
        (
            .in_data({
                         in_data[237],
                         in_data[89],
                         in_data[278],
                         in_data[506],
                         in_data[771],
                         in_data[209]
                    }),
            .out_data(lut_306_out)
        );

reg   lut_306_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_306_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_306_ff <= lut_306_out;
    end
end

assign out_data[306] = lut_306_ff;




// LUT : 307

wire lut_307_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100111010010000110101110001000001010101111100000101011100110000),
            .DEVICE(DEVICE)
        )
    i_lut_307
        (
            .in_data({
                         in_data[452],
                         in_data[536],
                         in_data[676],
                         in_data[431],
                         in_data[777],
                         in_data[555]
                    }),
            .out_data(lut_307_out)
        );

reg   lut_307_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_307_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_307_ff <= lut_307_out;
    end
end

assign out_data[307] = lut_307_ff;




// LUT : 308

wire lut_308_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100001101000100100100100000000011001000101001111010110000010011),
            .DEVICE(DEVICE)
        )
    i_lut_308
        (
            .in_data({
                         in_data[217],
                         in_data[358],
                         in_data[446],
                         in_data[562],
                         in_data[270],
                         in_data[123]
                    }),
            .out_data(lut_308_out)
        );

reg   lut_308_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_308_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_308_ff <= lut_308_out;
    end
end

assign out_data[308] = lut_308_ff;




// LUT : 309

wire lut_309_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110011011111110001101110111111110100000011100101011101010111111),
            .DEVICE(DEVICE)
        )
    i_lut_309
        (
            .in_data({
                         in_data[409],
                         in_data[207],
                         in_data[287],
                         in_data[227],
                         in_data[114],
                         in_data[239]
                    }),
            .out_data(lut_309_out)
        );

reg   lut_309_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_309_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_309_ff <= lut_309_out;
    end
end

assign out_data[309] = lut_309_ff;




// LUT : 310

wire lut_310_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010110100110100010000010000001000011111010111110111011101111),
            .DEVICE(DEVICE)
        )
    i_lut_310
        (
            .in_data({
                         in_data[722],
                         in_data[193],
                         in_data[208],
                         in_data[42],
                         in_data[691],
                         in_data[422]
                    }),
            .out_data(lut_310_out)
        );

reg   lut_310_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_310_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_310_ff <= lut_310_out;
    end
end

assign out_data[310] = lut_310_ff;




// LUT : 311

wire lut_311_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010111010101100000000001101110010100110001011001001100001111),
            .DEVICE(DEVICE)
        )
    i_lut_311
        (
            .in_data({
                         in_data[651],
                         in_data[268],
                         in_data[685],
                         in_data[746],
                         in_data[566],
                         in_data[440]
                    }),
            .out_data(lut_311_out)
        );

reg   lut_311_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_311_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_311_ff <= lut_311_out;
    end
end

assign out_data[311] = lut_311_ff;




// LUT : 312

wire lut_312_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100010101111110101101100000001010000010100001110000001011000),
            .DEVICE(DEVICE)
        )
    i_lut_312
        (
            .in_data({
                         in_data[360],
                         in_data[336],
                         in_data[101],
                         in_data[656],
                         in_data[780],
                         in_data[94]
                    }),
            .out_data(lut_312_out)
        );

reg   lut_312_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_312_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_312_ff <= lut_312_out;
    end
end

assign out_data[312] = lut_312_ff;




// LUT : 313

wire lut_313_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010111010110000101110100111010111011110101111101000110000000),
            .DEVICE(DEVICE)
        )
    i_lut_313
        (
            .in_data({
                         in_data[453],
                         in_data[558],
                         in_data[252],
                         in_data[385],
                         in_data[546],
                         in_data[76]
                    }),
            .out_data(lut_313_out)
        );

reg   lut_313_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_313_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_313_ff <= lut_313_out;
    end
end

assign out_data[313] = lut_313_ff;




// LUT : 314

wire lut_314_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010011111000011000110000000110001001101100101111010110110100),
            .DEVICE(DEVICE)
        )
    i_lut_314
        (
            .in_data({
                         in_data[504],
                         in_data[726],
                         in_data[66],
                         in_data[172],
                         in_data[550],
                         in_data[510]
                    }),
            .out_data(lut_314_out)
        );

reg   lut_314_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_314_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_314_ff <= lut_314_out;
    end
end

assign out_data[314] = lut_314_ff;




// LUT : 315

wire lut_315_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001010000100000001111000000100011101101100000100111101100011),
            .DEVICE(DEVICE)
        )
    i_lut_315
        (
            .in_data({
                         in_data[773],
                         in_data[621],
                         in_data[586],
                         in_data[69],
                         in_data[282],
                         in_data[265]
                    }),
            .out_data(lut_315_out)
        );

reg   lut_315_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_315_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_315_ff <= lut_315_out;
    end
end

assign out_data[315] = lut_315_ff;




// LUT : 316

wire lut_316_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000100000110001011111111011101110001000100010111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_316
        (
            .in_data({
                         in_data[734],
                         in_data[156],
                         in_data[299],
                         in_data[486],
                         in_data[118],
                         in_data[326]
                    }),
            .out_data(lut_316_out)
        );

reg   lut_316_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_316_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_316_ff <= lut_316_out;
    end
end

assign out_data[316] = lut_316_ff;




// LUT : 317

wire lut_317_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100011100101011110001001000000100111001101100011110100111000),
            .DEVICE(DEVICE)
        )
    i_lut_317
        (
            .in_data({
                         in_data[142],
                         in_data[88],
                         in_data[383],
                         in_data[333],
                         in_data[748],
                         in_data[604]
                    }),
            .out_data(lut_317_out)
        );

reg   lut_317_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_317_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_317_ff <= lut_317_out;
    end
end

assign out_data[317] = lut_317_ff;




// LUT : 318

wire lut_318_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001000011110011010010101100111000000011101001000010110011101),
            .DEVICE(DEVICE)
        )
    i_lut_318
        (
            .in_data({
                         in_data[571],
                         in_data[744],
                         in_data[548],
                         in_data[697],
                         in_data[618],
                         in_data[703]
                    }),
            .out_data(lut_318_out)
        );

reg   lut_318_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_318_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_318_ff <= lut_318_out;
    end
end

assign out_data[318] = lut_318_ff;




// LUT : 319

wire lut_319_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100100101100111111101101100100111101001010001111100110001000),
            .DEVICE(DEVICE)
        )
    i_lut_319
        (
            .in_data({
                         in_data[12],
                         in_data[508],
                         in_data[574],
                         in_data[692],
                         in_data[747],
                         in_data[11]
                    }),
            .out_data(lut_319_out)
        );

reg   lut_319_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_319_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_319_ff <= lut_319_out;
    end
end

assign out_data[319] = lut_319_ff;




// LUT : 320

wire lut_320_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101001101001010101001110111001011000001101110010000110100111110),
            .DEVICE(DEVICE)
        )
    i_lut_320
        (
            .in_data({
                         in_data[567],
                         in_data[553],
                         in_data[32],
                         in_data[110],
                         in_data[355],
                         in_data[166]
                    }),
            .out_data(lut_320_out)
        );

reg   lut_320_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_320_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_320_ff <= lut_320_out;
    end
end

assign out_data[320] = lut_320_ff;




// LUT : 321

wire lut_321_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000010000000100010001000000010101010001000001000000010000001),
            .DEVICE(DEVICE)
        )
    i_lut_321
        (
            .in_data({
                         in_data[176],
                         in_data[180],
                         in_data[528],
                         in_data[663],
                         in_data[624],
                         in_data[92]
                    }),
            .out_data(lut_321_out)
        );

reg   lut_321_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_321_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_321_ff <= lut_321_out;
    end
end

assign out_data[321] = lut_321_ff;




// LUT : 322

wire lut_322_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010111011101111011100001011111000010101000001100010010001101),
            .DEVICE(DEVICE)
        )
    i_lut_322
        (
            .in_data({
                         in_data[345],
                         in_data[414],
                         in_data[471],
                         in_data[151],
                         in_data[285],
                         in_data[25]
                    }),
            .out_data(lut_322_out)
        );

reg   lut_322_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_322_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_322_ff <= lut_322_out;
    end
end

assign out_data[322] = lut_322_ff;




// LUT : 323

wire lut_323_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100101010001000000101001000000001000111000000111111111100000111),
            .DEVICE(DEVICE)
        )
    i_lut_323
        (
            .in_data({
                         in_data[466],
                         in_data[485],
                         in_data[342],
                         in_data[233],
                         in_data[334],
                         in_data[687]
                    }),
            .out_data(lut_323_out)
        );

reg   lut_323_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_323_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_323_ff <= lut_323_out;
    end
end

assign out_data[323] = lut_323_ff;




// LUT : 324

wire lut_324_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010101000100111111111111111100111001000100110101010111011111),
            .DEVICE(DEVICE)
        )
    i_lut_324
        (
            .in_data({
                         in_data[328],
                         in_data[413],
                         in_data[186],
                         in_data[210],
                         in_data[584],
                         in_data[293]
                    }),
            .out_data(lut_324_out)
        );

reg   lut_324_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_324_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_324_ff <= lut_324_out;
    end
end

assign out_data[324] = lut_324_ff;




// LUT : 325

wire lut_325_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010011011111001001111100010111110000001101010111101110100100),
            .DEVICE(DEVICE)
        )
    i_lut_325
        (
            .in_data({
                         in_data[753],
                         in_data[313],
                         in_data[384],
                         in_data[645],
                         in_data[731],
                         in_data[614]
                    }),
            .out_data(lut_325_out)
        );

reg   lut_325_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_325_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_325_ff <= lut_325_out;
    end
end

assign out_data[325] = lut_325_ff;




// LUT : 326

wire lut_326_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100001101010011111011011100010010111010110111001001100010000),
            .DEVICE(DEVICE)
        )
    i_lut_326
        (
            .in_data({
                         in_data[769],
                         in_data[82],
                         in_data[41],
                         in_data[23],
                         in_data[218],
                         in_data[236]
                    }),
            .out_data(lut_326_out)
        );

reg   lut_326_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_326_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_326_ff <= lut_326_out;
    end
end

assign out_data[326] = lut_326_ff;




// LUT : 327

wire lut_327_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011110100000111110010001100110111100101001101101011110110001111),
            .DEVICE(DEVICE)
        )
    i_lut_327
        (
            .in_data({
                         in_data[640],
                         in_data[14],
                         in_data[420],
                         in_data[192],
                         in_data[484],
                         in_data[9]
                    }),
            .out_data(lut_327_out)
        );

reg   lut_327_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_327_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_327_ff <= lut_327_out;
    end
end

assign out_data[327] = lut_327_ff;




// LUT : 328

wire lut_328_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000101011100011100111001101011101010100100000001011011011010),
            .DEVICE(DEVICE)
        )
    i_lut_328
        (
            .in_data({
                         in_data[526],
                         in_data[671],
                         in_data[124],
                         in_data[447],
                         in_data[759],
                         in_data[93]
                    }),
            .out_data(lut_328_out)
        );

reg   lut_328_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_328_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_328_ff <= lut_328_out;
    end
end

assign out_data[328] = lut_328_ff;




// LUT : 329

wire lut_329_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100111111011101111111101110010101011010111111001101101111100),
            .DEVICE(DEVICE)
        )
    i_lut_329
        (
            .in_data({
                         in_data[382],
                         in_data[261],
                         in_data[195],
                         in_data[13],
                         in_data[179],
                         in_data[712]
                    }),
            .out_data(lut_329_out)
        );

reg   lut_329_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_329_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_329_ff <= lut_329_out;
    end
end

assign out_data[329] = lut_329_ff;




// LUT : 330

wire lut_330_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110101010000101100011111000111110000000001001111101100011111),
            .DEVICE(DEVICE)
        )
    i_lut_330
        (
            .in_data({
                         in_data[106],
                         in_data[455],
                         in_data[601],
                         in_data[147],
                         in_data[509],
                         in_data[520]
                    }),
            .out_data(lut_330_out)
        );

reg   lut_330_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_330_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_330_ff <= lut_330_out;
    end
end

assign out_data[330] = lut_330_ff;




// LUT : 331

wire lut_331_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001011010010000100101101001110100010111110101011001011110011),
            .DEVICE(DEVICE)
        )
    i_lut_331
        (
            .in_data({
                         in_data[636],
                         in_data[605],
                         in_data[439],
                         in_data[444],
                         in_data[398],
                         in_data[525]
                    }),
            .out_data(lut_331_out)
        );

reg   lut_331_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_331_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_331_ff <= lut_331_out;
    end
end

assign out_data[331] = lut_331_ff;




// LUT : 332

wire lut_332_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101011001110111001101101100000001011100010111010101101111111),
            .DEVICE(DEVICE)
        )
    i_lut_332
        (
            .in_data({
                         in_data[719],
                         in_data[74],
                         in_data[73],
                         in_data[609],
                         in_data[595],
                         in_data[450]
                    }),
            .out_data(lut_332_out)
        );

reg   lut_332_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_332_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_332_ff <= lut_332_out;
    end
end

assign out_data[332] = lut_332_ff;




// LUT : 333

wire lut_333_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001001010110111011010101101000001100110101011111100001011010101),
            .DEVICE(DEVICE)
        )
    i_lut_333
        (
            .in_data({
                         in_data[259],
                         in_data[122],
                         in_data[778],
                         in_data[369],
                         in_data[776],
                         in_data[146]
                    }),
            .out_data(lut_333_out)
        );

reg   lut_333_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_333_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_333_ff <= lut_333_out;
    end
end

assign out_data[333] = lut_333_ff;




// LUT : 334

wire lut_334_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100101110100111010100000111101110111111011000110010111111101),
            .DEVICE(DEVICE)
        )
    i_lut_334
        (
            .in_data({
                         in_data[353],
                         in_data[34],
                         in_data[701],
                         in_data[113],
                         in_data[26],
                         in_data[538]
                    }),
            .out_data(lut_334_out)
        );

reg   lut_334_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_334_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_334_ff <= lut_334_out;
    end
end

assign out_data[334] = lut_334_ff;




// LUT : 335

wire lut_335_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000100011101110000110101001110011001110001000000101001000100101),
            .DEVICE(DEVICE)
        )
    i_lut_335
        (
            .in_data({
                         in_data[655],
                         in_data[330],
                         in_data[620],
                         in_data[63],
                         in_data[544],
                         in_data[308]
                    }),
            .out_data(lut_335_out)
        );

reg   lut_335_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_335_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_335_ff <= lut_335_out;
    end
end

assign out_data[335] = lut_335_ff;




// LUT : 336

wire lut_336_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101100001100101111000000001010100001111010101010000011010101),
            .DEVICE(DEVICE)
        )
    i_lut_336
        (
            .in_data({
                         in_data[433],
                         in_data[763],
                         in_data[738],
                         in_data[304],
                         in_data[593],
                         in_data[153]
                    }),
            .out_data(lut_336_out)
        );

reg   lut_336_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_336_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_336_ff <= lut_336_out;
    end
end

assign out_data[336] = lut_336_ff;




// LUT : 337

wire lut_337_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100111101111101011011010000001001110011111111111100011111101),
            .DEVICE(DEVICE)
        )
    i_lut_337
        (
            .in_data({
                         in_data[626],
                         in_data[432],
                         in_data[17],
                         in_data[411],
                         in_data[44],
                         in_data[202]
                    }),
            .out_data(lut_337_out)
        );

reg   lut_337_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_337_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_337_ff <= lut_337_out;
    end
end

assign out_data[337] = lut_337_ff;




// LUT : 338

wire lut_338_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111011101111001010000100110010101111011111110100111110111100),
            .DEVICE(DEVICE)
        )
    i_lut_338
        (
            .in_data({
                         in_data[684],
                         in_data[181],
                         in_data[535],
                         in_data[38],
                         in_data[598],
                         in_data[325]
                    }),
            .out_data(lut_338_out)
        );

reg   lut_338_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_338_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_338_ff <= lut_338_out;
    end
end

assign out_data[338] = lut_338_ff;




// LUT : 339

wire lut_339_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101001111110110100001001000000001011011010100110011110111111111),
            .DEVICE(DEVICE)
        )
    i_lut_339
        (
            .in_data({
                         in_data[137],
                         in_data[650],
                         in_data[599],
                         in_data[589],
                         in_data[770],
                         in_data[511]
                    }),
            .out_data(lut_339_out)
        );

reg   lut_339_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_339_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_339_ff <= lut_339_out;
    end
end

assign out_data[339] = lut_339_ff;




// LUT : 340

wire lut_340_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101111011100111101001001010011110001100011011100110001011111),
            .DEVICE(DEVICE)
        )
    i_lut_340
        (
            .in_data({
                         in_data[628],
                         in_data[649],
                         in_data[664],
                         in_data[752],
                         in_data[395],
                         in_data[633]
                    }),
            .out_data(lut_340_out)
        );

reg   lut_340_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_340_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_340_ff <= lut_340_out;
    end
end

assign out_data[340] = lut_340_ff;




// LUT : 341

wire lut_341_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001011111000110011101111111111111111111111111011111010101000),
            .DEVICE(DEVICE)
        )
    i_lut_341
        (
            .in_data({
                         in_data[250],
                         in_data[160],
                         in_data[472],
                         in_data[515],
                         in_data[573],
                         in_data[578]
                    }),
            .out_data(lut_341_out)
        );

reg   lut_341_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_341_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_341_ff <= lut_341_out;
    end
end

assign out_data[341] = lut_341_ff;




// LUT : 342

wire lut_342_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100011101011111101101011000110111010101011111111111010101110101),
            .DEVICE(DEVICE)
        )
    i_lut_342
        (
            .in_data({
                         in_data[152],
                         in_data[373],
                         in_data[603],
                         in_data[721],
                         in_data[606],
                         in_data[463]
                    }),
            .out_data(lut_342_out)
        );

reg   lut_342_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_342_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_342_ff <= lut_342_out;
    end
end

assign out_data[342] = lut_342_ff;




// LUT : 343

wire lut_343_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110011010100111011000110101010100000001100101001001100111110110),
            .DEVICE(DEVICE)
        )
    i_lut_343
        (
            .in_data({
                         in_data[499],
                         in_data[662],
                         in_data[754],
                         in_data[419],
                         in_data[500],
                         in_data[563]
                    }),
            .out_data(lut_343_out)
        );

reg   lut_343_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_343_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_343_ff <= lut_343_out;
    end
end

assign out_data[343] = lut_343_ff;




// LUT : 344

wire lut_344_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001100100111100011000001010110100100010111111000100100010101),
            .DEVICE(DEVICE)
        )
    i_lut_344
        (
            .in_data({
                         in_data[232],
                         in_data[575],
                         in_data[51],
                         in_data[407],
                         in_data[518],
                         in_data[762]
                    }),
            .out_data(lut_344_out)
        );

reg   lut_344_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_344_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_344_ff <= lut_344_out;
    end
end

assign out_data[344] = lut_344_ff;




// LUT : 345

wire lut_345_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000011000110110100111011010100011001011011011101011000000010),
            .DEVICE(DEVICE)
        )
    i_lut_345
        (
            .in_data({
                         in_data[613],
                         in_data[706],
                         in_data[112],
                         in_data[311],
                         in_data[430],
                         in_data[693]
                    }),
            .out_data(lut_345_out)
        );

reg   lut_345_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_345_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_345_ff <= lut_345_out;
    end
end

assign out_data[345] = lut_345_ff;




// LUT : 346

wire lut_346_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001100000010010011011000001110011111000000100110110101100011),
            .DEVICE(DEVICE)
        )
    i_lut_346
        (
            .in_data({
                         in_data[681],
                         in_data[482],
                         in_data[699],
                         in_data[495],
                         in_data[612],
                         in_data[581]
                    }),
            .out_data(lut_346_out)
        );

reg   lut_346_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_346_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_346_ff <= lut_346_out;
    end
end

assign out_data[346] = lut_346_ff;




// LUT : 347

wire lut_347_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011110010111001011101110100010001010001111010111011100100110),
            .DEVICE(DEVICE)
        )
    i_lut_347
        (
            .in_data({
                         in_data[381],
                         in_data[46],
                         in_data[322],
                         in_data[460],
                         in_data[729],
                         in_data[657]
                    }),
            .out_data(lut_347_out)
        );

reg   lut_347_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_347_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_347_ff <= lut_347_out;
    end
end

assign out_data[347] = lut_347_ff;




// LUT : 348

wire lut_348_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011111001010111001001010010100010100111011110110100110111110),
            .DEVICE(DEVICE)
        )
    i_lut_348
        (
            .in_data({
                         in_data[675],
                         in_data[203],
                         in_data[20],
                         in_data[62],
                         in_data[229],
                         in_data[674]
                    }),
            .out_data(lut_348_out)
        );

reg   lut_348_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_348_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_348_ff <= lut_348_out;
    end
end

assign out_data[348] = lut_348_ff;




// LUT : 349

wire lut_349_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010101100111000000010000001111110101001000110011010010001110),
            .DEVICE(DEVICE)
        )
    i_lut_349
        (
            .in_data({
                         in_data[677],
                         in_data[512],
                         in_data[324],
                         in_data[37],
                         in_data[412],
                         in_data[481]
                    }),
            .out_data(lut_349_out)
        );

reg   lut_349_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_349_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_349_ff <= lut_349_out;
    end
end

assign out_data[349] = lut_349_ff;




// LUT : 350

wire lut_350_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100010000011110110110100011000001100011011100001000100000001),
            .DEVICE(DEVICE)
        )
    i_lut_350
        (
            .in_data({
                         in_data[255],
                         in_data[61],
                         in_data[545],
                         in_data[461],
                         in_data[277],
                         in_data[221]
                    }),
            .out_data(lut_350_out)
        );

reg   lut_350_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_350_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_350_ff <= lut_350_out;
    end
end

assign out_data[350] = lut_350_ff;




// LUT : 351

wire lut_351_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010010100000101100101000010000100111000100100101110100001000),
            .DEVICE(DEVICE)
        )
    i_lut_351
        (
            .in_data({
                         in_data[591],
                         in_data[19],
                         in_data[387],
                         in_data[349],
                         in_data[1],
                         in_data[351]
                    }),
            .out_data(lut_351_out)
        );

reg   lut_351_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_351_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_351_ff <= lut_351_out;
    end
end

assign out_data[351] = lut_351_ff;




// LUT : 352

wire lut_352_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010011010100101100001101100100010001101111101010110100010100100),
            .DEVICE(DEVICE)
        )
    i_lut_352
        (
            .in_data({
                         in_data[178],
                         in_data[28],
                         in_data[368],
                         in_data[300],
                         in_data[139],
                         in_data[80]
                    }),
            .out_data(lut_352_out)
        );

reg   lut_352_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_352_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_352_ff <= lut_352_out;
    end
end

assign out_data[352] = lut_352_ff;




// LUT : 353

wire lut_353_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101101000111011110110110011010011011011101011011101111110011),
            .DEVICE(DEVICE)
        )
    i_lut_353
        (
            .in_data({
                         in_data[272],
                         in_data[402],
                         in_data[710],
                         in_data[540],
                         in_data[128],
                         in_data[264]
                    }),
            .out_data(lut_353_out)
        );

reg   lut_353_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_353_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_353_ff <= lut_353_out;
    end
end

assign out_data[353] = lut_353_ff;




// LUT : 354

wire lut_354_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100111110001110101011011110110000101100001110101000010001100),
            .DEVICE(DEVICE)
        )
    i_lut_354
        (
            .in_data({
                         in_data[281],
                         in_data[241],
                         in_data[258],
                         in_data[266],
                         in_data[196],
                         in_data[52]
                    }),
            .out_data(lut_354_out)
        );

reg   lut_354_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_354_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_354_ff <= lut_354_out;
    end
end

assign out_data[354] = lut_354_ff;




// LUT : 355

wire lut_355_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101111111101010011110011111110110001110001001010100111100111),
            .DEVICE(DEVICE)
        )
    i_lut_355
        (
            .in_data({
                         in_data[145],
                         in_data[290],
                         in_data[5],
                         in_data[428],
                         in_data[537],
                         in_data[492]
                    }),
            .out_data(lut_355_out)
        );

reg   lut_355_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_355_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_355_ff <= lut_355_out;
    end
end

assign out_data[355] = lut_355_ff;




// LUT : 356

wire lut_356_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000000001111000010101100100001100110111001000000101010001100),
            .DEVICE(DEVICE)
        )
    i_lut_356
        (
            .in_data({
                         in_data[119],
                         in_data[404],
                         in_data[223],
                         in_data[27],
                         in_data[6],
                         in_data[117]
                    }),
            .out_data(lut_356_out)
        );

reg   lut_356_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_356_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_356_ff <= lut_356_out;
    end
end

assign out_data[356] = lut_356_ff;




// LUT : 357

wire lut_357_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100011101001100110011010100101011010010010101101010010100101010),
            .DEVICE(DEVICE)
        )
    i_lut_357
        (
            .in_data({
                         in_data[523],
                         in_data[83],
                         in_data[457],
                         in_data[58],
                         in_data[376],
                         in_data[253]
                    }),
            .out_data(lut_357_out)
        );

reg   lut_357_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_357_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_357_ff <= lut_357_out;
    end
end

assign out_data[357] = lut_357_ff;




// LUT : 358

wire lut_358_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000111010100100111000000000101101101011110011010101101101011),
            .DEVICE(DEVICE)
        )
    i_lut_358
        (
            .in_data({
                         in_data[163],
                         in_data[554],
                         in_data[109],
                         in_data[7],
                         in_data[531],
                         in_data[449]
                    }),
            .out_data(lut_358_out)
        );

reg   lut_358_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_358_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_358_ff <= lut_358_out;
    end
end

assign out_data[358] = lut_358_ff;




// LUT : 359

wire lut_359_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111111000000111110111001010001100110011000110111110001000101),
            .DEVICE(DEVICE)
        )
    i_lut_359
        (
            .in_data({
                         in_data[339],
                         in_data[48],
                         in_data[54],
                         in_data[617],
                         in_data[646],
                         in_data[86]
                    }),
            .out_data(lut_359_out)
        );

reg   lut_359_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_359_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_359_ff <= lut_359_out;
    end
end

assign out_data[359] = lut_359_ff;




// LUT : 360

wire lut_360_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110001001000010101011011000111100000001001001111101011111100),
            .DEVICE(DEVICE)
        )
    i_lut_360
        (
            .in_data({
                         in_data[517],
                         in_data[425],
                         in_data[458],
                         in_data[36],
                         in_data[775],
                         in_data[696]
                    }),
            .out_data(lut_360_out)
        );

reg   lut_360_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_360_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_360_ff <= lut_360_out;
    end
end

assign out_data[360] = lut_360_ff;




// LUT : 361

wire lut_361_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111110110100010001000111000111101001111111011101111011110111),
            .DEVICE(DEVICE)
        )
    i_lut_361
        (
            .in_data({
                         in_data[427],
                         in_data[585],
                         in_data[50],
                         in_data[779],
                         in_data[724],
                         in_data[582]
                    }),
            .out_data(lut_361_out)
        );

reg   lut_361_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_361_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_361_ff <= lut_361_out;
    end
end

assign out_data[361] = lut_361_ff;




// LUT : 362

wire lut_362_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000100010001110011000001100101110011001000101111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_362
        (
            .in_data({
                         in_data[451],
                         in_data[317],
                         in_data[228],
                         in_data[435],
                         in_data[718],
                         in_data[256]
                    }),
            .out_data(lut_362_out)
        );

reg   lut_362_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_362_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_362_ff <= lut_362_out;
    end
end

assign out_data[362] = lut_362_ff;




// LUT : 363

wire lut_363_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111101100010000000000000100101100011110011100000000010110111),
            .DEVICE(DEVICE)
        )
    i_lut_363
        (
            .in_data({
                         in_data[442],
                         in_data[115],
                         in_data[415],
                         in_data[214],
                         in_data[246],
                         in_data[204]
                    }),
            .out_data(lut_363_out)
        );

reg   lut_363_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_363_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_363_ff <= lut_363_out;
    end
end

assign out_data[363] = lut_363_ff;




// LUT : 364

wire lut_364_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110000000110111100010011011101100011010001011110110000000001010),
            .DEVICE(DEVICE)
        )
    i_lut_364
        (
            .in_data({
                         in_data[488],
                         in_data[619],
                         in_data[338],
                         in_data[332],
                         in_data[388],
                         in_data[379]
                    }),
            .out_data(lut_364_out)
        );

reg   lut_364_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_364_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_364_ff <= lut_364_out;
    end
end

assign out_data[364] = lut_364_ff;




// LUT : 365

wire lut_365_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100101101101100110110000000010011010010010000100101010110011),
            .DEVICE(DEVICE)
        )
    i_lut_365
        (
            .in_data({
                         in_data[743],
                         in_data[104],
                         in_data[138],
                         in_data[372],
                         in_data[170],
                         in_data[354]
                    }),
            .out_data(lut_365_out)
        );

reg   lut_365_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_365_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_365_ff <= lut_365_out;
    end
end

assign out_data[365] = lut_365_ff;




// LUT : 366

wire lut_366_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011110111010110111001000011001010111010001111110100101000001101),
            .DEVICE(DEVICE)
        )
    i_lut_366
        (
            .in_data({
                         in_data[77],
                         in_data[105],
                         in_data[198],
                         in_data[67],
                         in_data[723],
                         in_data[647]
                    }),
            .out_data(lut_366_out)
        );

reg   lut_366_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_366_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_366_ff <= lut_366_out;
    end
end

assign out_data[366] = lut_366_ff;




// LUT : 367

wire lut_367_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100111011111000001111000010000010110111000101100111100100000),
            .DEVICE(DEVICE)
        )
    i_lut_367
        (
            .in_data({
                         in_data[288],
                         in_data[21],
                         in_data[527],
                         in_data[760],
                         in_data[594],
                         in_data[197]
                    }),
            .out_data(lut_367_out)
        );

reg   lut_367_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_367_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_367_ff <= lut_367_out;
    end
end

assign out_data[367] = lut_367_ff;




// LUT : 368

wire lut_368_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100101001110011100110001110100001111110111110001111000011110),
            .DEVICE(DEVICE)
        )
    i_lut_368
        (
            .in_data({
                         in_data[100],
                         in_data[749],
                         in_data[319],
                         in_data[49],
                         in_data[725],
                         in_data[296]
                    }),
            .out_data(lut_368_out)
        );

reg   lut_368_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_368_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_368_ff <= lut_368_out;
    end
end

assign out_data[368] = lut_368_ff;




// LUT : 369

wire lut_369_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010001010001000110000000011011100000011010000000101001110000),
            .DEVICE(DEVICE)
        )
    i_lut_369
        (
            .in_data({
                         in_data[426],
                         in_data[251],
                         in_data[745],
                         in_data[700],
                         in_data[758],
                         in_data[167]
                    }),
            .out_data(lut_369_out)
        );

reg   lut_369_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_369_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_369_ff <= lut_369_out;
    end
end

assign out_data[369] = lut_369_ff;




// LUT : 370

wire lut_370_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100110000101000100000101100110101111000011111100111101001111),
            .DEVICE(DEVICE)
        )
    i_lut_370
        (
            .in_data({
                         in_data[560],
                         in_data[271],
                         in_data[654],
                         in_data[549],
                         in_data[741],
                         in_data[519]
                    }),
            .out_data(lut_370_out)
        );

reg   lut_370_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_370_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_370_ff <= lut_370_out;
    end
end

assign out_data[370] = lut_370_ff;




// LUT : 371

wire lut_371_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011101111011100011001100001100001000000010100101101011111010),
            .DEVICE(DEVICE)
        )
    i_lut_371
        (
            .in_data({
                         in_data[740],
                         in_data[68],
                         in_data[361],
                         in_data[199],
                         in_data[580],
                         in_data[213]
                    }),
            .out_data(lut_371_out)
        );

reg   lut_371_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_371_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_371_ff <= lut_371_out;
    end
end

assign out_data[371] = lut_371_ff;




// LUT : 372

wire lut_372_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001111011111001101001011111110101111000010101011101100110111),
            .DEVICE(DEVICE)
        )
    i_lut_372
        (
            .in_data({
                         in_data[474],
                         in_data[183],
                         in_data[648],
                         in_data[344],
                         in_data[157],
                         in_data[177]
                    }),
            .out_data(lut_372_out)
        );

reg   lut_372_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_372_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_372_ff <= lut_372_out;
    end
end

assign out_data[372] = lut_372_ff;




// LUT : 373

wire lut_373_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100010001011000011011100111101000001110101010000000001000100),
            .DEVICE(DEVICE)
        )
    i_lut_373
        (
            .in_data({
                         in_data[689],
                         in_data[507],
                         in_data[742],
                         in_data[539],
                         in_data[10],
                         in_data[374]
                    }),
            .out_data(lut_373_out)
        );

reg   lut_373_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_373_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_373_ff <= lut_373_out;
    end
end

assign out_data[373] = lut_373_ff;




// LUT : 374

wire lut_374_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000101000101010101011101111101111100110101010111101010100010),
            .DEVICE(DEVICE)
        )
    i_lut_374
        (
            .in_data({
                         in_data[524],
                         in_data[362],
                         in_data[454],
                         in_data[348],
                         in_data[576],
                         in_data[18]
                    }),
            .out_data(lut_374_out)
        );

reg   lut_374_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_374_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_374_ff <= lut_374_out;
    end
end

assign out_data[374] = lut_374_ff;




// LUT : 375

wire lut_375_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101011000000110111110000000011111010000110111111101000010011),
            .DEVICE(DEVICE)
        )
    i_lut_375
        (
            .in_data({
                         in_data[371],
                         in_data[263],
                         in_data[136],
                         in_data[274],
                         in_data[347],
                         in_data[470]
                    }),
            .out_data(lut_375_out)
        );

reg   lut_375_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_375_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_375_ff <= lut_375_out;
    end
end

assign out_data[375] = lut_375_ff;




// LUT : 376

wire lut_376_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100010111010011111011111110101011111110111011101011100101110),
            .DEVICE(DEVICE)
        )
    i_lut_376
        (
            .in_data({
                         in_data[249],
                         in_data[561],
                         in_data[248],
                         in_data[456],
                         in_data[627],
                         in_data[225]
                    }),
            .out_data(lut_376_out)
        );

reg   lut_376_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_376_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_376_ff <= lut_376_out;
    end
end

assign out_data[376] = lut_376_ff;




// LUT : 377

wire lut_377_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111110100101100101000000101111100110001111011000110000000001),
            .DEVICE(DEVICE)
        )
    i_lut_377
        (
            .in_data({
                         in_data[15],
                         in_data[364],
                         in_data[212],
                         in_data[331],
                         in_data[55],
                         in_data[135]
                    }),
            .out_data(lut_377_out)
        );

reg   lut_377_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_377_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_377_ff <= lut_377_out;
    end
end

assign out_data[377] = lut_377_ff;




// LUT : 378

wire lut_378_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100100101110001001001101110001001100001110111000100001010101),
            .DEVICE(DEVICE)
        )
    i_lut_378
        (
            .in_data({
                         in_data[502],
                         in_data[565],
                         in_data[401],
                         in_data[188],
                         in_data[335],
                         in_data[498]
                    }),
            .out_data(lut_378_out)
        );

reg   lut_378_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_378_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_378_ff <= lut_378_out;
    end
end

assign out_data[378] = lut_378_ff;




// LUT : 379

wire lut_379_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000100000000000111110001000000000000111000000100110011000101101),
            .DEVICE(DEVICE)
        )
    i_lut_379
        (
            .in_data({
                         in_data[514],
                         in_data[634],
                         in_data[683],
                         in_data[162],
                         in_data[405],
                         in_data[559]
                    }),
            .out_data(lut_379_out)
        );

reg   lut_379_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_379_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_379_ff <= lut_379_out;
    end
end

assign out_data[379] = lut_379_ff;




// LUT : 380

wire lut_380_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110000000010100111000000000000000011000001011000000000000101),
            .DEVICE(DEVICE)
        )
    i_lut_380
        (
            .in_data({
                         in_data[120],
                         in_data[610],
                         in_data[478],
                         in_data[97],
                         in_data[185],
                         in_data[327]
                    }),
            .out_data(lut_380_out)
        );

reg   lut_380_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_380_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_380_ff <= lut_380_out;
    end
end

assign out_data[380] = lut_380_ff;




// LUT : 381

wire lut_381_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001000100010110010100111011101111101110100011011101011000111),
            .DEVICE(DEVICE)
        )
    i_lut_381
        (
            .in_data({
                         in_data[400],
                         in_data[24],
                         in_data[483],
                         in_data[33],
                         in_data[489],
                         in_data[702]
                    }),
            .out_data(lut_381_out)
        );

reg   lut_381_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_381_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_381_ff <= lut_381_out;
    end
end

assign out_data[381] = lut_381_ff;




// LUT : 382

wire lut_382_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000010011010101011011000100101000111011011000000000111001010),
            .DEVICE(DEVICE)
        )
    i_lut_382
        (
            .in_data({
                         in_data[238],
                         in_data[533],
                         in_data[698],
                         in_data[493],
                         in_data[4],
                         in_data[216]
                    }),
            .out_data(lut_382_out)
        );

reg   lut_382_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_382_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_382_ff <= lut_382_out;
    end
end

assign out_data[382] = lut_382_ff;




// LUT : 383

wire lut_383_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110010010101110001010100110110100100000001011100011011000101),
            .DEVICE(DEVICE)
        )
    i_lut_383
        (
            .in_data({
                         in_data[568],
                         in_data[494],
                         in_data[448],
                         in_data[389],
                         in_data[39],
                         in_data[244]
                    }),
            .out_data(lut_383_out)
        );

reg   lut_383_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_383_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_383_ff <= lut_383_out;
    end
end

assign out_data[383] = lut_383_ff;




// LUT : 384

wire lut_384_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111011011001010010010101011101101000100101101010001000101011),
            .DEVICE(DEVICE)
        )
    i_lut_384
        (
            .in_data({
                         in_data[730],
                         in_data[30],
                         in_data[564],
                         in_data[148],
                         in_data[301],
                         in_data[0]
                    }),
            .out_data(lut_384_out)
        );

reg   lut_384_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_384_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_384_ff <= lut_384_out;
    end
end

assign out_data[384] = lut_384_ff;




// LUT : 385

wire lut_385_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100001001111100101010001001101101010011010001110110010100111101),
            .DEVICE(DEVICE)
        )
    i_lut_385
        (
            .in_data({
                         in_data[226],
                         in_data[764],
                         in_data[149],
                         in_data[783],
                         in_data[781],
                         in_data[140]
                    }),
            .out_data(lut_385_out)
        );

reg   lut_385_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_385_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_385_ff <= lut_385_out;
    end
end

assign out_data[385] = lut_385_ff;




// LUT : 386

wire lut_386_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011100101010000111011001100000011010001011010110101001000101),
            .DEVICE(DEVICE)
        )
    i_lut_386
        (
            .in_data({
                         in_data[670],
                         in_data[359],
                         in_data[480],
                         in_data[280],
                         in_data[403],
                         in_data[768]
                    }),
            .out_data(lut_386_out)
        );

reg   lut_386_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_386_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_386_ff <= lut_386_out;
    end
end

assign out_data[386] = lut_386_ff;




// LUT : 387

wire lut_387_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010011110010011101110010011001110110100101000110001111000001000),
            .DEVICE(DEVICE)
        )
    i_lut_387
        (
            .in_data({
                         in_data[386],
                         in_data[184],
                         in_data[84],
                         in_data[245],
                         in_data[200],
                         in_data[739]
                    }),
            .out_data(lut_387_out)
        );

reg   lut_387_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_387_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_387_ff <= lut_387_out;
    end
end

assign out_data[387] = lut_387_ff;




// LUT : 388

wire lut_388_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100011111010000001101110000001000001011011000100011111110110),
            .DEVICE(DEVICE)
        )
    i_lut_388
        (
            .in_data({
                         in_data[468],
                         in_data[2],
                         in_data[211],
                         in_data[755],
                         in_data[732],
                         in_data[108]
                    }),
            .out_data(lut_388_out)
        );

reg   lut_388_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_388_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_388_ff <= lut_388_out;
    end
end

assign out_data[388] = lut_388_ff;




// LUT : 389

wire lut_389_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101011110001100100101101000011101100110000111111001110000011),
            .DEVICE(DEVICE)
        )
    i_lut_389
        (
            .in_data({
                         in_data[716],
                         in_data[590],
                         in_data[592],
                         in_data[394],
                         in_data[206],
                         in_data[174]
                    }),
            .out_data(lut_389_out)
        );

reg   lut_389_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_389_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_389_ff <= lut_389_out;
    end
end

assign out_data[389] = lut_389_ff;




// LUT : 390

wire lut_390_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010000111100110110010011100100011100100110011010000001000000),
            .DEVICE(DEVICE)
        )
    i_lut_390
        (
            .in_data({
                         in_data[634],
                         in_data[781],
                         in_data[437],
                         in_data[60],
                         in_data[475],
                         in_data[445]
                    }),
            .out_data(lut_390_out)
        );

reg   lut_390_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_390_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_390_ff <= lut_390_out;
    end
end

assign out_data[390] = lut_390_ff;




// LUT : 391

wire lut_391_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000110001010111111001011101011101010010000000000011000001010110),
            .DEVICE(DEVICE)
        )
    i_lut_391
        (
            .in_data({
                         in_data[518],
                         in_data[356],
                         in_data[0],
                         in_data[316],
                         in_data[21],
                         in_data[284]
                    }),
            .out_data(lut_391_out)
        );

reg   lut_391_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_391_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_391_ff <= lut_391_out;
    end
end

assign out_data[391] = lut_391_ff;




// LUT : 392

wire lut_392_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001111101110011100001011111111110010001111000110111011010111),
            .DEVICE(DEVICE)
        )
    i_lut_392
        (
            .in_data({
                         in_data[278],
                         in_data[45],
                         in_data[33],
                         in_data[595],
                         in_data[366],
                         in_data[552]
                    }),
            .out_data(lut_392_out)
        );

reg   lut_392_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_392_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_392_ff <= lut_392_out;
    end
end

assign out_data[392] = lut_392_ff;




// LUT : 393

wire lut_393_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000011010001100010001010001001101010010101111111101111001101),
            .DEVICE(DEVICE)
        )
    i_lut_393
        (
            .in_data({
                         in_data[590],
                         in_data[701],
                         in_data[5],
                         in_data[180],
                         in_data[714],
                         in_data[560]
                    }),
            .out_data(lut_393_out)
        );

reg   lut_393_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_393_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_393_ff <= lut_393_out;
    end
end

assign out_data[393] = lut_393_ff;




// LUT : 394

wire lut_394_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111001010001110011110011011010000001110101010110101100110110),
            .DEVICE(DEVICE)
        )
    i_lut_394
        (
            .in_data({
                         in_data[288],
                         in_data[503],
                         in_data[530],
                         in_data[359],
                         in_data[112],
                         in_data[734]
                    }),
            .out_data(lut_394_out)
        );

reg   lut_394_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_394_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_394_ff <= lut_394_out;
    end
end

assign out_data[394] = lut_394_ff;




// LUT : 395

wire lut_395_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110101000100111110111010101111110010010111110111110110000000100),
            .DEVICE(DEVICE)
        )
    i_lut_395
        (
            .in_data({
                         in_data[721],
                         in_data[227],
                         in_data[512],
                         in_data[588],
                         in_data[543],
                         in_data[674]
                    }),
            .out_data(lut_395_out)
        );

reg   lut_395_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_395_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_395_ff <= lut_395_out;
    end
end

assign out_data[395] = lut_395_ff;




// LUT : 396

wire lut_396_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101000100101001010000011001110110101101101111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_396
        (
            .in_data({
                         in_data[140],
                         in_data[103],
                         in_data[155],
                         in_data[237],
                         in_data[171],
                         in_data[174]
                    }),
            .out_data(lut_396_out)
        );

reg   lut_396_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_396_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_396_ff <= lut_396_out;
    end
end

assign out_data[396] = lut_396_ff;




// LUT : 397

wire lut_397_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111110011011111000011000111111111001000001100110100110010001100),
            .DEVICE(DEVICE)
        )
    i_lut_397
        (
            .in_data({
                         in_data[344],
                         in_data[347],
                         in_data[447],
                         in_data[461],
                         in_data[28],
                         in_data[91]
                    }),
            .out_data(lut_397_out)
        );

reg   lut_397_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_397_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_397_ff <= lut_397_out;
    end
end

assign out_data[397] = lut_397_ff;




// LUT : 398

wire lut_398_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010110011111111101111101111110010000111001111111111101010111100),
            .DEVICE(DEVICE)
        )
    i_lut_398
        (
            .in_data({
                         in_data[492],
                         in_data[746],
                         in_data[651],
                         in_data[220],
                         in_data[282],
                         in_data[352]
                    }),
            .out_data(lut_398_out)
        );

reg   lut_398_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_398_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_398_ff <= lut_398_out;
    end
end

assign out_data[398] = lut_398_ff;




// LUT : 399

wire lut_399_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000001000100000000000110011101100110011001100110010),
            .DEVICE(DEVICE)
        )
    i_lut_399
        (
            .in_data({
                         in_data[520],
                         in_data[272],
                         in_data[259],
                         in_data[686],
                         in_data[738],
                         in_data[273]
                    }),
            .out_data(lut_399_out)
        );

reg   lut_399_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_399_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_399_ff <= lut_399_out;
    end
end

assign out_data[399] = lut_399_ff;




// LUT : 400

wire lut_400_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001011111110000001111100101011100000001001100000111110100001),
            .DEVICE(DEVICE)
        )
    i_lut_400
        (
            .in_data({
                         in_data[717],
                         in_data[42],
                         in_data[453],
                         in_data[185],
                         in_data[10],
                         in_data[110]
                    }),
            .out_data(lut_400_out)
        );

reg   lut_400_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_400_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_400_ff <= lut_400_out;
    end
end

assign out_data[400] = lut_400_ff;




// LUT : 401

wire lut_401_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000001010000101100000001000100000000110101010110000110000111),
            .DEVICE(DEVICE)
        )
    i_lut_401
        (
            .in_data({
                         in_data[154],
                         in_data[657],
                         in_data[631],
                         in_data[113],
                         in_data[331],
                         in_data[228]
                    }),
            .out_data(lut_401_out)
        );

reg   lut_401_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_401_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_401_ff <= lut_401_out;
    end
end

assign out_data[401] = lut_401_ff;




// LUT : 402

wire lut_402_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000101010000011001101101000110101000111100000000111000110111),
            .DEVICE(DEVICE)
        )
    i_lut_402
        (
            .in_data({
                         in_data[574],
                         in_data[609],
                         in_data[187],
                         in_data[770],
                         in_data[51],
                         in_data[204]
                    }),
            .out_data(lut_402_out)
        );

reg   lut_402_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_402_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_402_ff <= lut_402_out;
    end
end

assign out_data[402] = lut_402_ff;




// LUT : 403

wire lut_403_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110011111011101010010101111011001100001111111010101101001110010),
            .DEVICE(DEVICE)
        )
    i_lut_403
        (
            .in_data({
                         in_data[209],
                         in_data[41],
                         in_data[747],
                         in_data[441],
                         in_data[765],
                         in_data[478]
                    }),
            .out_data(lut_403_out)
        );

reg   lut_403_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_403_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_403_ff <= lut_403_out;
    end
end

assign out_data[403] = lut_403_ff;




// LUT : 404

wire lut_404_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011110100111011011001011101011111010000101000110010101000111010),
            .DEVICE(DEVICE)
        )
    i_lut_404
        (
            .in_data({
                         in_data[371],
                         in_data[16],
                         in_data[567],
                         in_data[731],
                         in_data[539],
                         in_data[100]
                    }),
            .out_data(lut_404_out)
        );

reg   lut_404_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_404_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_404_ff <= lut_404_out;
    end
end

assign out_data[404] = lut_404_ff;




// LUT : 405

wire lut_405_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000000111110101100010101000110010011111101100001101110111111),
            .DEVICE(DEVICE)
        )
    i_lut_405
        (
            .in_data({
                         in_data[732],
                         in_data[604],
                         in_data[446],
                         in_data[568],
                         in_data[368],
                         in_data[696]
                    }),
            .out_data(lut_405_out)
        );

reg   lut_405_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_405_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_405_ff <= lut_405_out;
    end
end

assign out_data[405] = lut_405_ff;




// LUT : 406

wire lut_406_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010000110010111000101011000011111110000011011101011001000111),
            .DEVICE(DEVICE)
        )
    i_lut_406
        (
            .in_data({
                         in_data[58],
                         in_data[689],
                         in_data[725],
                         in_data[691],
                         in_data[349],
                         in_data[654]
                    }),
            .out_data(lut_406_out)
        );

reg   lut_406_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_406_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_406_ff <= lut_406_out;
    end
end

assign out_data[406] = lut_406_ff;




// LUT : 407

wire lut_407_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100001001110101000100011101101110001011001111110011100100000),
            .DEVICE(DEVICE)
        )
    i_lut_407
        (
            .in_data({
                         in_data[418],
                         in_data[666],
                         in_data[728],
                         in_data[15],
                         in_data[358],
                         in_data[53]
                    }),
            .out_data(lut_407_out)
        );

reg   lut_407_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_407_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_407_ff <= lut_407_out;
    end
end

assign out_data[407] = lut_407_ff;




// LUT : 408

wire lut_408_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010010010001111000101000100110111000101110111000100000111111),
            .DEVICE(DEVICE)
        )
    i_lut_408
        (
            .in_data({
                         in_data[381],
                         in_data[501],
                         in_data[306],
                         in_data[429],
                         in_data[274],
                         in_data[671]
                    }),
            .out_data(lut_408_out)
        );

reg   lut_408_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_408_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_408_ff <= lut_408_out;
    end
end

assign out_data[408] = lut_408_ff;




// LUT : 409

wire lut_409_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110111011111011100010000000000011001000001011101110010000100000),
            .DEVICE(DEVICE)
        )
    i_lut_409
        (
            .in_data({
                         in_data[542],
                         in_data[678],
                         in_data[493],
                         in_data[267],
                         in_data[223],
                         in_data[462]
                    }),
            .out_data(lut_409_out)
        );

reg   lut_409_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_409_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_409_ff <= lut_409_out;
    end
end

assign out_data[409] = lut_409_ff;




// LUT : 410

wire lut_410_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111110111111101111001111110001111100111111000011010010111101),
            .DEVICE(DEVICE)
        )
    i_lut_410
        (
            .in_data({
                         in_data[291],
                         in_data[287],
                         in_data[385],
                         in_data[771],
                         in_data[777],
                         in_data[383]
                    }),
            .out_data(lut_410_out)
        );

reg   lut_410_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_410_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_410_ff <= lut_410_out;
    end
end

assign out_data[410] = lut_410_ff;




// LUT : 411

wire lut_411_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011110001101001101111010100101011101001100010111000101110100),
            .DEVICE(DEVICE)
        )
    i_lut_411
        (
            .in_data({
                         in_data[338],
                         in_data[162],
                         in_data[555],
                         in_data[242],
                         in_data[225],
                         in_data[29]
                    }),
            .out_data(lut_411_out)
        );

reg   lut_411_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_411_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_411_ff <= lut_411_out;
    end
end

assign out_data[411] = lut_411_ff;




// LUT : 412

wire lut_412_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011110010100110100001100010011001111101111001110110001001100000),
            .DEVICE(DEVICE)
        )
    i_lut_412
        (
            .in_data({
                         in_data[334],
                         in_data[415],
                         in_data[136],
                         in_data[144],
                         in_data[135],
                         in_data[69]
                    }),
            .out_data(lut_412_out)
        );

reg   lut_412_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_412_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_412_ff <= lut_412_out;
    end
end

assign out_data[412] = lut_412_ff;




// LUT : 413

wire lut_413_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001100101100011110110001010101110000111010110011001100100100010),
            .DEVICE(DEVICE)
        )
    i_lut_413
        (
            .in_data({
                         in_data[217],
                         in_data[733],
                         in_data[7],
                         in_data[336],
                         in_data[40],
                         in_data[362]
                    }),
            .out_data(lut_413_out)
        );

reg   lut_413_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_413_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_413_ff <= lut_413_out;
    end
end

assign out_data[413] = lut_413_ff;




// LUT : 414

wire lut_414_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001001101110010000110101001001110010010011000010000011001100),
            .DEVICE(DEVICE)
        )
    i_lut_414
        (
            .in_data({
                         in_data[584],
                         in_data[427],
                         in_data[193],
                         in_data[759],
                         in_data[212],
                         in_data[663]
                    }),
            .out_data(lut_414_out)
        );

reg   lut_414_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_414_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_414_ff <= lut_414_out;
    end
end

assign out_data[414] = lut_414_ff;




// LUT : 415

wire lut_415_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011011001111010101100011110000111111110001100100111010100110),
            .DEVICE(DEVICE)
        )
    i_lut_415
        (
            .in_data({
                         in_data[55],
                         in_data[684],
                         in_data[495],
                         in_data[54],
                         in_data[6],
                         in_data[249]
                    }),
            .out_data(lut_415_out)
        );

reg   lut_415_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_415_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_415_ff <= lut_415_out;
    end
end

assign out_data[415] = lut_415_ff;




// LUT : 416

wire lut_416_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001001100000000000010000000001000000001000000000000001000000101),
            .DEVICE(DEVICE)
        )
    i_lut_416
        (
            .in_data({
                         in_data[471],
                         in_data[64],
                         in_data[467],
                         in_data[457],
                         in_data[326],
                         in_data[36]
                    }),
            .out_data(lut_416_out)
        );

reg   lut_416_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_416_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_416_ff <= lut_416_out;
    end
end

assign out_data[416] = lut_416_ff;




// LUT : 417

wire lut_417_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010000111101000100001101000101100100001101010100010000010000),
            .DEVICE(DEVICE)
        )
    i_lut_417
        (
            .in_data({
                         in_data[121],
                         in_data[353],
                         in_data[425],
                         in_data[350],
                         in_data[750],
                         in_data[544]
                    }),
            .out_data(lut_417_out)
        );

reg   lut_417_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_417_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_417_ff <= lut_417_out;
    end
end

assign out_data[417] = lut_417_ff;




// LUT : 418

wire lut_418_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100101001100011011101011010000001101100010000100000001000110),
            .DEVICE(DEVICE)
        )
    i_lut_418
        (
            .in_data({
                         in_data[409],
                         in_data[585],
                         in_data[66],
                         in_data[498],
                         in_data[22],
                         in_data[693]
                    }),
            .out_data(lut_418_out)
        );

reg   lut_418_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_418_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_418_ff <= lut_418_out;
    end
end

assign out_data[418] = lut_418_ff;




// LUT : 419

wire lut_419_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111001100110000001110000001111111101111101100110011101111),
            .DEVICE(DEVICE)
        )
    i_lut_419
        (
            .in_data({
                         in_data[569],
                         in_data[563],
                         in_data[258],
                         in_data[201],
                         in_data[687],
                         in_data[215]
                    }),
            .out_data(lut_419_out)
        );

reg   lut_419_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_419_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_419_ff <= lut_419_out;
    end
end

assign out_data[419] = lut_419_ff;




// LUT : 420

wire lut_420_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110111000001110111111111111111111101000101111111010011111010),
            .DEVICE(DEVICE)
        )
    i_lut_420
        (
            .in_data({
                         in_data[536],
                         in_data[198],
                         in_data[188],
                         in_data[608],
                         in_data[514],
                         in_data[147]
                    }),
            .out_data(lut_420_out)
        );

reg   lut_420_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_420_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_420_ff <= lut_420_out;
    end
end

assign out_data[420] = lut_420_ff;




// LUT : 421

wire lut_421_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010001110100000011111000111011000000111000001111111101011000),
            .DEVICE(DEVICE)
        )
    i_lut_421
        (
            .in_data({
                         in_data[145],
                         in_data[489],
                         in_data[294],
                         in_data[422],
                         in_data[321],
                         in_data[148]
                    }),
            .out_data(lut_421_out)
        );

reg   lut_421_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_421_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_421_ff <= lut_421_out;
    end
end

assign out_data[421] = lut_421_ff;




// LUT : 422

wire lut_422_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111011100000111100001001000010100110101001100110110011000111),
            .DEVICE(DEVICE)
        )
    i_lut_422
        (
            .in_data({
                         in_data[76],
                         in_data[405],
                         in_data[434],
                         in_data[618],
                         in_data[165],
                         in_data[395]
                    }),
            .out_data(lut_422_out)
        );

reg   lut_422_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_422_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_422_ff <= lut_422_out;
    end
end

assign out_data[422] = lut_422_ff;




// LUT : 423

wire lut_423_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100110110011100001110011101100110010111110001011111100110000),
            .DEVICE(DEVICE)
        )
    i_lut_423
        (
            .in_data({
                         in_data[531],
                         in_data[472],
                         in_data[301],
                         in_data[458],
                         in_data[256],
                         in_data[176]
                    }),
            .out_data(lut_423_out)
        );

reg   lut_423_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_423_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_423_ff <= lut_423_out;
    end
end

assign out_data[423] = lut_423_ff;




// LUT : 424

wire lut_424_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111000100011011000011010000111000111111100111000101111110011),
            .DEVICE(DEVICE)
        )
    i_lut_424
        (
            .in_data({
                         in_data[276],
                         in_data[236],
                         in_data[311],
                         in_data[77],
                         in_data[428],
                         in_data[160]
                    }),
            .out_data(lut_424_out)
        );

reg   lut_424_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_424_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_424_ff <= lut_424_out;
    end
end

assign out_data[424] = lut_424_ff;




// LUT : 425

wire lut_425_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111110101010101111110011101000011111101111110111111101111111),
            .DEVICE(DEVICE)
        )
    i_lut_425
        (
            .in_data({
                         in_data[516],
                         in_data[407],
                         in_data[715],
                         in_data[255],
                         in_data[443],
                         in_data[414]
                    }),
            .out_data(lut_425_out)
        );

reg   lut_425_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_425_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_425_ff <= lut_425_out;
    end
end

assign out_data[425] = lut_425_ff;




// LUT : 426

wire lut_426_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110000010001110001010001110110000100001101011111010000110101100),
            .DEVICE(DEVICE)
        )
    i_lut_426
        (
            .in_data({
                         in_data[75],
                         in_data[372],
                         in_data[402],
                         in_data[742],
                         in_data[424],
                         in_data[124]
                    }),
            .out_data(lut_426_out)
        );

reg   lut_426_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_426_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_426_ff <= lut_426_out;
    end
end

assign out_data[426] = lut_426_ff;




// LUT : 427

wire lut_427_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011110011001110000110110101000101100100101000101010110010011),
            .DEVICE(DEVICE)
        )
    i_lut_427
        (
            .in_data({
                         in_data[80],
                         in_data[554],
                         in_data[111],
                         in_data[599],
                         in_data[707],
                         in_data[122]
                    }),
            .out_data(lut_427_out)
        );

reg   lut_427_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_427_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_427_ff <= lut_427_out;
    end
end

assign out_data[427] = lut_427_ff;




// LUT : 428

wire lut_428_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100001001000101100111111111101001110111011100111011001110001000),
            .DEVICE(DEVICE)
        )
    i_lut_428
        (
            .in_data({
                         in_data[169],
                         in_data[736],
                         in_data[292],
                         in_data[632],
                         in_data[783],
                         in_data[626]
                    }),
            .out_data(lut_428_out)
        );

reg   lut_428_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_428_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_428_ff <= lut_428_out;
    end
end

assign out_data[428] = lut_428_ff;




// LUT : 429

wire lut_429_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110000101110010001000000000011011111010001000101110111001100),
            .DEVICE(DEVICE)
        )
    i_lut_429
        (
            .in_data({
                         in_data[213],
                         in_data[35],
                         in_data[440],
                         in_data[581],
                         in_data[384],
                         in_data[150]
                    }),
            .out_data(lut_429_out)
        );

reg   lut_429_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_429_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_429_ff <= lut_429_out;
    end
end

assign out_data[429] = lut_429_ff;




// LUT : 430

wire lut_430_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111001110111101011010011110101000000110101000000000101010101),
            .DEVICE(DEVICE)
        )
    i_lut_430
        (
            .in_data({
                         in_data[720],
                         in_data[466],
                         in_data[751],
                         in_data[444],
                         in_data[183],
                         in_data[95]
                    }),
            .out_data(lut_430_out)
        );

reg   lut_430_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_430_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_430_ff <= lut_430_out;
    end
end

assign out_data[430] = lut_430_ff;




// LUT : 431

wire lut_431_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110000101010100101100101011010111110110101101101111000110110),
            .DEVICE(DEVICE)
        )
    i_lut_431
        (
            .in_data({
                         in_data[98],
                         in_data[591],
                         in_data[374],
                         in_data[191],
                         in_data[723],
                         in_data[309]
                    }),
            .out_data(lut_431_out)
        );

reg   lut_431_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_431_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_431_ff <= lut_431_out;
    end
end

assign out_data[431] = lut_431_ff;




// LUT : 432

wire lut_432_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111100000011110111101000000010111111110111101000100010000001),
            .DEVICE(DEVICE)
        )
    i_lut_432
        (
            .in_data({
                         in_data[342],
                         in_data[729],
                         in_data[647],
                         in_data[605],
                         in_data[59],
                         in_data[547]
                    }),
            .out_data(lut_432_out)
        );

reg   lut_432_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_432_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_432_ff <= lut_432_out;
    end
end

assign out_data[432] = lut_432_ff;




// LUT : 433

wire lut_433_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101000110110000000100001100011111111101110111111101011111010),
            .DEVICE(DEVICE)
        )
    i_lut_433
        (
            .in_data({
                         in_data[318],
                         in_data[580],
                         in_data[433],
                         in_data[635],
                         in_data[119],
                         in_data[583]
                    }),
            .out_data(lut_433_out)
        );

reg   lut_433_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_433_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_433_ff <= lut_433_out;
    end
end

assign out_data[433] = lut_433_ff;




// LUT : 434

wire lut_434_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010101000101001001010100010100000101000001001100110100000100),
            .DEVICE(DEVICE)
        )
    i_lut_434
        (
            .in_data({
                         in_data[206],
                         in_data[189],
                         in_data[650],
                         in_data[137],
                         in_data[577],
                         in_data[345]
                    }),
            .out_data(lut_434_out)
        );

reg   lut_434_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_434_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_434_ff <= lut_434_out;
    end
end

assign out_data[434] = lut_434_ff;




// LUT : 435

wire lut_435_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000001011000111101011100101000111100101110101110111000010101),
            .DEVICE(DEVICE)
        )
    i_lut_435
        (
            .in_data({
                         in_data[613],
                         in_data[640],
                         in_data[365],
                         in_data[172],
                         in_data[92],
                         in_data[194]
                    }),
            .out_data(lut_435_out)
        );

reg   lut_435_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_435_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_435_ff <= lut_435_out;
    end
end

assign out_data[435] = lut_435_ff;




// LUT : 436

wire lut_436_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100111100001101110100111000000011000001001010010010000011000000),
            .DEVICE(DEVICE)
        )
    i_lut_436
        (
            .in_data({
                         in_data[315],
                         in_data[570],
                         in_data[252],
                         in_data[247],
                         in_data[11],
                         in_data[339]
                    }),
            .out_data(lut_436_out)
        );

reg   lut_436_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_436_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_436_ff <= lut_436_out;
    end
end

assign out_data[436] = lut_436_ff;




// LUT : 437

wire lut_437_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111011111110111111101111111101111111011111110),
            .DEVICE(DEVICE)
        )
    i_lut_437
        (
            .in_data({
                         in_data[178],
                         in_data[628],
                         in_data[602],
                         in_data[411],
                         in_data[302],
                         in_data[578]
                    }),
            .out_data(lut_437_out)
        );

reg   lut_437_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_437_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_437_ff <= lut_437_out;
    end
end

assign out_data[437] = lut_437_ff;




// LUT : 438

wire lut_438_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101100000101011000000000010100101000001000011100001010000011),
            .DEVICE(DEVICE)
        )
    i_lut_438
        (
            .in_data({
                         in_data[261],
                         in_data[603],
                         in_data[62],
                         in_data[184],
                         in_data[233],
                         in_data[744]
                    }),
            .out_data(lut_438_out)
        );

reg   lut_438_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_438_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_438_ff <= lut_438_out;
    end
end

assign out_data[438] = lut_438_ff;




// LUT : 439

wire lut_439_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001000001010101011101111111111010101010000000011001100000001),
            .DEVICE(DEVICE)
        )
    i_lut_439
        (
            .in_data({
                         in_data[1],
                         in_data[50],
                         in_data[639],
                         in_data[438],
                         in_data[768],
                         in_data[576]
                    }),
            .out_data(lut_439_out)
        );

reg   lut_439_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_439_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_439_ff <= lut_439_out;
    end
end

assign out_data[439] = lut_439_ff;




// LUT : 440

wire lut_440_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110111101110101101011000100011001010101110111010010001011101100),
            .DEVICE(DEVICE)
        )
    i_lut_440
        (
            .in_data({
                         in_data[549],
                         in_data[297],
                         in_data[523],
                         in_data[575],
                         in_data[661],
                         in_data[17]
                    }),
            .out_data(lut_440_out)
        );

reg   lut_440_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_440_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_440_ff <= lut_440_out;
    end
end

assign out_data[440] = lut_440_ff;




// LUT : 441

wire lut_441_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111001101101001111110101011110111110010001101110001011101010),
            .DEVICE(DEVICE)
        )
    i_lut_441
        (
            .in_data({
                         in_data[99],
                         in_data[665],
                         in_data[521],
                         in_data[699],
                         in_data[592],
                         in_data[323]
                    }),
            .out_data(lut_441_out)
        );

reg   lut_441_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_441_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_441_ff <= lut_441_out;
    end
end

assign out_data[441] = lut_441_ff;




// LUT : 442

wire lut_442_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110101100110111010101110010101100100100000011000100010000011001),
            .DEVICE(DEVICE)
        )
    i_lut_442
        (
            .in_data({
                         in_data[329],
                         in_data[659],
                         in_data[545],
                         in_data[586],
                         in_data[34],
                         in_data[293]
                    }),
            .out_data(lut_442_out)
        );

reg   lut_442_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_442_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_442_ff <= lut_442_out;
    end
end

assign out_data[442] = lut_442_ff;




// LUT : 443

wire lut_443_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000000100000001000000100010001110000000001101111100011101110),
            .DEVICE(DEVICE)
        )
    i_lut_443
        (
            .in_data({
                         in_data[120],
                         in_data[151],
                         in_data[67],
                         in_data[44],
                         in_data[214],
                         in_data[566]
                    }),
            .out_data(lut_443_out)
        );

reg   lut_443_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_443_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_443_ff <= lut_443_out;
    end
end

assign out_data[443] = lut_443_ff;




// LUT : 444

wire lut_444_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111000010100000010001110100000001010111101001110111010111001),
            .DEVICE(DEVICE)
        )
    i_lut_444
        (
            .in_data({
                         in_data[504],
                         in_data[668],
                         in_data[515],
                         in_data[295],
                         in_data[27],
                         in_data[56]
                    }),
            .out_data(lut_444_out)
        );

reg   lut_444_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_444_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_444_ff <= lut_444_out;
    end
end

assign out_data[444] = lut_444_ff;




// LUT : 445

wire lut_445_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001100000010000010111110110011101011011010000000001101101010),
            .DEVICE(DEVICE)
        )
    i_lut_445
        (
            .in_data({
                         in_data[465],
                         in_data[662],
                         in_data[317],
                         in_data[506],
                         in_data[14],
                         in_data[389]
                    }),
            .out_data(lut_445_out)
        );

reg   lut_445_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_445_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_445_ff <= lut_445_out;
    end
end

assign out_data[445] = lut_445_ff;




// LUT : 446

wire lut_446_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000111010010101010000101000011101101111010010110000011001000),
            .DEVICE(DEVICE)
        )
    i_lut_446
        (
            .in_data({
                         in_data[403],
                         in_data[623],
                         in_data[745],
                         in_data[752],
                         in_data[420],
                         in_data[398]
                    }),
            .out_data(lut_446_out)
        );

reg   lut_446_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_446_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_446_ff <= lut_446_out;
    end
end

assign out_data[446] = lut_446_ff;




// LUT : 447

wire lut_447_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101100110011011011110100001111111111111011111111100010111000),
            .DEVICE(DEVICE)
        )
    i_lut_447
        (
            .in_data({
                         in_data[199],
                         in_data[128],
                         in_data[638],
                         in_data[219],
                         in_data[508],
                         in_data[431]
                    }),
            .out_data(lut_447_out)
        );

reg   lut_447_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_447_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_447_ff <= lut_447_out;
    end
end

assign out_data[447] = lut_447_ff;




// LUT : 448

wire lut_448_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010000000110001101110110011101000110000110001011101111111111),
            .DEVICE(DEVICE)
        )
    i_lut_448
        (
            .in_data({
                         in_data[529],
                         in_data[248],
                         in_data[179],
                         in_data[679],
                         in_data[129],
                         in_data[81]
                    }),
            .out_data(lut_448_out)
        );

reg   lut_448_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_448_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_448_ff <= lut_448_out;
    end
end

assign out_data[448] = lut_448_ff;




// LUT : 449

wire lut_449_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001001010100000110000100000000000100010100100000101011110010000),
            .DEVICE(DEVICE)
        )
    i_lut_449
        (
            .in_data({
                         in_data[455],
                         in_data[63],
                         in_data[488],
                         in_data[540],
                         in_data[413],
                         in_data[669]
                    }),
            .out_data(lut_449_out)
        );

reg   lut_449_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_449_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_449_ff <= lut_449_out;
    end
end

assign out_data[449] = lut_449_ff;




// LUT : 450

wire lut_450_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010101100101111010111001010010100001100111110011101000000100),
            .DEVICE(DEVICE)
        )
    i_lut_450
        (
            .in_data({
                         in_data[268],
                         in_data[304],
                         in_data[97],
                         in_data[26],
                         in_data[724],
                         in_data[43]
                    }),
            .out_data(lut_450_out)
        );

reg   lut_450_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_450_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_450_ff <= lut_450_out;
    end
end

assign out_data[450] = lut_450_ff;




// LUT : 451

wire lut_451_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001111011011000111001000010101011101101100011100110111011100110),
            .DEVICE(DEVICE)
        )
    i_lut_451
        (
            .in_data({
                         in_data[764],
                         in_data[727],
                         in_data[210],
                         in_data[386],
                         in_data[587],
                         in_data[460]
                    }),
            .out_data(lut_451_out)
        );

reg   lut_451_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_451_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_451_ff <= lut_451_out;
    end
end

assign out_data[451] = lut_451_ff;




// LUT : 452

wire lut_452_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010111111111010111010001101111001101100111110101111101011111),
            .DEVICE(DEVICE)
        )
    i_lut_452
        (
            .in_data({
                         in_data[468],
                         in_data[341],
                         in_data[553],
                         in_data[133],
                         in_data[325],
                         in_data[207]
                    }),
            .out_data(lut_452_out)
        );

reg   lut_452_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_452_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_452_ff <= lut_452_out;
    end
end

assign out_data[452] = lut_452_ff;




// LUT : 453

wire lut_453_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111001111010010011011011000000111110011100011001001100010110000),
            .DEVICE(DEVICE)
        )
    i_lut_453
        (
            .in_data({
                         in_data[82],
                         in_data[704],
                         in_data[68],
                         in_data[483],
                         in_data[627],
                         in_data[528]
                    }),
            .out_data(lut_453_out)
        );

reg   lut_453_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_453_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_453_ff <= lut_453_out;
    end
end

assign out_data[453] = lut_453_ff;




// LUT : 454

wire lut_454_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011011001010100011101100010011110101011100000010101011011100),
            .DEVICE(DEVICE)
        )
    i_lut_454
        (
            .in_data({
                         in_data[675],
                         in_data[216],
                         in_data[226],
                         in_data[401],
                         in_data[633],
                         in_data[335]
                    }),
            .out_data(lut_454_out)
        );

reg   lut_454_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_454_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_454_ff <= lut_454_out;
    end
end

assign out_data[454] = lut_454_ff;




// LUT : 455

wire lut_455_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000011111100111101110111110001110101111100001111011101000100),
            .DEVICE(DEVICE)
        )
    i_lut_455
        (
            .in_data({
                         in_data[522],
                         in_data[509],
                         in_data[312],
                         in_data[367],
                         in_data[308],
                         in_data[396]
                    }),
            .out_data(lut_455_out)
        );

reg   lut_455_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_455_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_455_ff <= lut_455_out;
    end
end

assign out_data[455] = lut_455_ff;




// LUT : 456

wire lut_456_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110111110010101000101101111110000000011011000010100011000100),
            .DEVICE(DEVICE)
        )
    i_lut_456
        (
            .in_data({
                         in_data[83],
                         in_data[410],
                         in_data[619],
                         in_data[181],
                         in_data[582],
                         in_data[281]
                    }),
            .out_data(lut_456_out)
        );

reg   lut_456_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_456_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_456_ff <= lut_456_out;
    end
end

assign out_data[456] = lut_456_ff;




// LUT : 457

wire lut_457_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111111000111100111011100111110001100001011001001110001011111),
            .DEVICE(DEVICE)
        )
    i_lut_457
        (
            .in_data({
                         in_data[322],
                         in_data[454],
                         in_data[426],
                         in_data[23],
                         in_data[221],
                         in_data[146]
                    }),
            .out_data(lut_457_out)
        );

reg   lut_457_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_457_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_457_ff <= lut_457_out;
    end
end

assign out_data[457] = lut_457_ff;




// LUT : 458

wire lut_458_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001011110110110001010111110100010101111101011111000110011001),
            .DEVICE(DEVICE)
        )
    i_lut_458
        (
            .in_data({
                         in_data[388],
                         in_data[57],
                         in_data[125],
                         in_data[534],
                         in_data[749],
                         in_data[2]
                    }),
            .out_data(lut_458_out)
        );

reg   lut_458_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_458_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_458_ff <= lut_458_out;
    end
end

assign out_data[458] = lut_458_ff;




// LUT : 459

wire lut_459_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000011100111001001011011000001001010111010000010010110100100),
            .DEVICE(DEVICE)
        )
    i_lut_459
        (
            .in_data({
                         in_data[391],
                         in_data[104],
                         in_data[269],
                         in_data[557],
                         in_data[205],
                         in_data[361]
                    }),
            .out_data(lut_459_out)
        );

reg   lut_459_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_459_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_459_ff <= lut_459_out;
    end
end

assign out_data[459] = lut_459_ff;




// LUT : 460

wire lut_460_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101001011011000010000101000101001000010010100000100011110101),
            .DEVICE(DEVICE)
        )
    i_lut_460
        (
            .in_data({
                         in_data[442],
                         in_data[157],
                         in_data[369],
                         in_data[156],
                         in_data[8],
                         in_data[392]
                    }),
            .out_data(lut_460_out)
        );

reg   lut_460_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_460_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_460_ff <= lut_460_out;
    end
end

assign out_data[460] = lut_460_ff;




// LUT : 461

wire lut_461_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110000100101000001010010010101111001001011100110100001100110111),
            .DEVICE(DEVICE)
        )
    i_lut_461
        (
            .in_data({
                         in_data[25],
                         in_data[115],
                         in_data[118],
                         in_data[589],
                         in_data[13],
                         in_data[562]
                    }),
            .out_data(lut_461_out)
        );

reg   lut_461_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_461_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_461_ff <= lut_461_out;
    end
end

assign out_data[461] = lut_461_ff;




// LUT : 462

wire lut_462_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100111011101110110110011101111101101110111111110011111110111),
            .DEVICE(DEVICE)
        )
    i_lut_462
        (
            .in_data({
                         in_data[307],
                         in_data[624],
                         in_data[319],
                         in_data[406],
                         in_data[480],
                         in_data[170]
                    }),
            .out_data(lut_462_out)
        );

reg   lut_462_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_462_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_462_ff <= lut_462_out;
    end
end

assign out_data[462] = lut_462_ff;




// LUT : 463

wire lut_463_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111101011101011101101100010100110111010001011110111110100000),
            .DEVICE(DEVICE)
        )
    i_lut_463
        (
            .in_data({
                         in_data[527],
                         in_data[132],
                         in_data[285],
                         in_data[251],
                         in_data[271],
                         in_data[450]
                    }),
            .out_data(lut_463_out)
        );

reg   lut_463_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_463_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_463_ff <= lut_463_out;
    end
end

assign out_data[463] = lut_463_ff;




// LUT : 464

wire lut_464_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111100100111100110010011111101101110000111000000011001111110),
            .DEVICE(DEVICE)
        )
    i_lut_464
        (
            .in_data({
                         in_data[629],
                         in_data[476],
                         in_data[298],
                         in_data[756],
                         in_data[594],
                         in_data[449]
                    }),
            .out_data(lut_464_out)
        );

reg   lut_464_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_464_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_464_ff <= lut_464_out;
    end
end

assign out_data[464] = lut_464_ff;




// LUT : 465

wire lut_465_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111101101110010111001100000010101001110001001000010101111110),
            .DEVICE(DEVICE)
        )
    i_lut_465
        (
            .in_data({
                         in_data[743],
                         in_data[253],
                         in_data[676],
                         in_data[484],
                         in_data[673],
                         in_data[46]
                    }),
            .out_data(lut_465_out)
        );

reg   lut_465_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_465_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_465_ff <= lut_465_out;
    end
end

assign out_data[465] = lut_465_ff;




// LUT : 466

wire lut_466_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101011000000111000010000010111011000000000001111000111100101),
            .DEVICE(DEVICE)
        )
    i_lut_466
        (
            .in_data({
                         in_data[463],
                         in_data[564],
                         in_data[257],
                         in_data[558],
                         in_data[517],
                         in_data[72]
                    }),
            .out_data(lut_466_out)
        );

reg   lut_466_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_466_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_466_ff <= lut_466_out;
    end
end

assign out_data[466] = lut_466_ff;




// LUT : 467

wire lut_467_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000111100010100110001011110000110011100101110001111011011110),
            .DEVICE(DEVICE)
        )
    i_lut_467
        (
            .in_data({
                         in_data[645],
                         in_data[737],
                         in_data[494],
                         in_data[93],
                         in_data[716],
                         in_data[741]
                    }),
            .out_data(lut_467_out)
        );

reg   lut_467_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_467_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_467_ff <= lut_467_out;
    end
end

assign out_data[467] = lut_467_ff;




// LUT : 468

wire lut_468_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000000000010100000000101000010010000111111101010000011110010),
            .DEVICE(DEVICE)
        )
    i_lut_468
        (
            .in_data({
                         in_data[740],
                         in_data[464],
                         in_data[203],
                         in_data[532],
                         in_data[290],
                         in_data[606]
                    }),
            .out_data(lut_468_out)
        );

reg   lut_468_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_468_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_468_ff <= lut_468_out;
    end
end

assign out_data[468] = lut_468_ff;




// LUT : 469

wire lut_469_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110011111111011111011111111000000010000000110010011010100111),
            .DEVICE(DEVICE)
        )
    i_lut_469
        (
            .in_data({
                         in_data[333],
                         in_data[435],
                         in_data[546],
                         in_data[652],
                         in_data[231],
                         in_data[755]
                    }),
            .out_data(lut_469_out)
        );

reg   lut_469_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_469_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_469_ff <= lut_469_out;
    end
end

assign out_data[469] = lut_469_ff;




// LUT : 470

wire lut_470_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111101010010111011111010100001100000111010000011010100111000),
            .DEVICE(DEVICE)
        )
    i_lut_470
        (
            .in_data({
                         in_data[234],
                         in_data[419],
                         in_data[763],
                         in_data[175],
                         in_data[131],
                         in_data[561]
                    }),
            .out_data(lut_470_out)
        );

reg   lut_470_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_470_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_470_ff <= lut_470_out;
    end
end

assign out_data[470] = lut_470_ff;




// LUT : 471

wire lut_471_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110001100111000111010011011000001101011101000111101111111111),
            .DEVICE(DEVICE)
        )
    i_lut_471
        (
            .in_data({
                         in_data[758],
                         in_data[351],
                         in_data[712],
                         in_data[706],
                         in_data[757],
                         in_data[238]
                    }),
            .out_data(lut_471_out)
        );

reg   lut_471_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_471_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_471_ff <= lut_471_out;
    end
end

assign out_data[471] = lut_471_ff;




// LUT : 472

wire lut_472_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110000101010111100111010011100000101000001011110101100111101),
            .DEVICE(DEVICE)
        )
    i_lut_472
        (
            .in_data({
                         in_data[642],
                         in_data[486],
                         in_data[102],
                         in_data[126],
                         in_data[664],
                         in_data[138]
                    }),
            .out_data(lut_472_out)
        );

reg   lut_472_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_472_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_472_ff <= lut_472_out;
    end
end

assign out_data[472] = lut_472_ff;




// LUT : 473

wire lut_473_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100010011111111011000001111111010101011111111001111001010011),
            .DEVICE(DEVICE)
        )
    i_lut_473
        (
            .in_data({
                         in_data[208],
                         in_data[596],
                         in_data[616],
                         in_data[116],
                         in_data[511],
                         in_data[346]
                    }),
            .out_data(lut_473_out)
        );

reg   lut_473_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_473_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_473_ff <= lut_473_out;
    end
end

assign out_data[473] = lut_473_ff;




// LUT : 474

wire lut_474_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001111101101010110100000001111111010010111000000011011100001),
            .DEVICE(DEVICE)
        )
    i_lut_474
        (
            .in_data({
                         in_data[481],
                         in_data[614],
                         in_data[718],
                         in_data[622],
                         in_data[767],
                         in_data[86]
                    }),
            .out_data(lut_474_out)
        );

reg   lut_474_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_474_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_474_ff <= lut_474_out;
    end
end

assign out_data[474] = lut_474_ff;




// LUT : 475

wire lut_475_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101011110110010010000010111111010011101011101110000111100000),
            .DEVICE(DEVICE)
        )
    i_lut_475
        (
            .in_data({
                         in_data[314],
                         in_data[108],
                         in_data[280],
                         in_data[142],
                         in_data[593],
                         in_data[513]
                    }),
            .out_data(lut_475_out)
        );

reg   lut_475_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_475_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_475_ff <= lut_475_out;
    end
end

assign out_data[475] = lut_475_ff;




// LUT : 476

wire lut_476_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111110111001001101101110011111101101111100100010111001100101011),
            .DEVICE(DEVICE)
        )
    i_lut_476
        (
            .in_data({
                         in_data[762],
                         in_data[615],
                         in_data[601],
                         in_data[692],
                         in_data[377],
                         in_data[761]
                    }),
            .out_data(lut_476_out)
        );

reg   lut_476_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_476_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_476_ff <= lut_476_out;
    end
end

assign out_data[476] = lut_476_ff;




// LUT : 477

wire lut_477_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111010110000001010010101010110111100010000110000111010001111),
            .DEVICE(DEVICE)
        )
    i_lut_477
        (
            .in_data({
                         in_data[730],
                         in_data[130],
                         in_data[173],
                         in_data[360],
                         in_data[690],
                         in_data[357]
                    }),
            .out_data(lut_477_out)
        );

reg   lut_477_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_477_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_477_ff <= lut_477_out;
    end
end

assign out_data[477] = lut_477_ff;




// LUT : 478

wire lut_478_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101011011100000001010000110001111010111110110011101010010010),
            .DEVICE(DEVICE)
        )
    i_lut_478
        (
            .in_data({
                         in_data[680],
                         in_data[695],
                         in_data[697],
                         in_data[12],
                         in_data[65],
                         in_data[196]
                    }),
            .out_data(lut_478_out)
        );

reg   lut_478_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_478_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_478_ff <= lut_478_out;
    end
end

assign out_data[478] = lut_478_ff;




// LUT : 479

wire lut_479_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000000100110001110010000011001110111011110101111000110110110),
            .DEVICE(DEVICE)
        )
    i_lut_479
        (
            .in_data({
                         in_data[393],
                         in_data[327],
                         in_data[330],
                         in_data[773],
                         in_data[134],
                         in_data[775]
                    }),
            .out_data(lut_479_out)
        );

reg   lut_479_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_479_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_479_ff <= lut_479_out;
    end
end

assign out_data[479] = lut_479_ff;




// LUT : 480

wire lut_480_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100010001011011110100111010000011111000001100101110000000100),
            .DEVICE(DEVICE)
        )
    i_lut_480
        (
            .in_data({
                         in_data[182],
                         in_data[222],
                         in_data[143],
                         in_data[753],
                         in_data[19],
                         in_data[477]
                    }),
            .out_data(lut_480_out)
        );

reg   lut_480_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_480_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_480_ff <= lut_480_out;
    end
end

assign out_data[480] = lut_480_ff;




// LUT : 481

wire lut_481_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100011110101000000101101010111101000001011110110010011110011110),
            .DEVICE(DEVICE)
        )
    i_lut_481
        (
            .in_data({
                         in_data[343],
                         in_data[735],
                         in_data[766],
                         in_data[32],
                         in_data[470],
                         in_data[778]
                    }),
            .out_data(lut_481_out)
        );

reg   lut_481_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_481_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_481_ff <= lut_481_out;
    end
end

assign out_data[481] = lut_481_ff;




// LUT : 482

wire lut_482_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010011101001001000101110011000011100110110001111111111101000),
            .DEVICE(DEVICE)
        )
    i_lut_482
        (
            .in_data({
                         in_data[535],
                         in_data[262],
                         in_data[340],
                         in_data[439],
                         in_data[620],
                         in_data[682]
                    }),
            .out_data(lut_482_out)
        );

reg   lut_482_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_482_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_482_ff <= lut_482_out;
    end
end

assign out_data[482] = lut_482_ff;




// LUT : 483

wire lut_483_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101001001100010110010000000101110011110011000101011111010111111),
            .DEVICE(DEVICE)
        )
    i_lut_483
        (
            .in_data({
                         in_data[127],
                         in_data[47],
                         in_data[378],
                         in_data[655],
                         in_data[260],
                         in_data[289]
                    }),
            .out_data(lut_483_out)
        );

reg   lut_483_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_483_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_483_ff <= lut_483_out;
    end
end

assign out_data[483] = lut_483_ff;




// LUT : 484

wire lut_484_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011010101111101111100010010011010000010000010001110000110001111),
            .DEVICE(DEVICE)
        )
    i_lut_484
        (
            .in_data({
                         in_data[355],
                         in_data[702],
                         in_data[79],
                         in_data[726],
                         in_data[611],
                         in_data[452]
                    }),
            .out_data(lut_484_out)
        );

reg   lut_484_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_484_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_484_ff <= lut_484_out;
    end
end

assign out_data[484] = lut_484_ff;




// LUT : 485

wire lut_485_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000110110001000011111100010101001000111111011000001011010011),
            .DEVICE(DEVICE)
        )
    i_lut_485
        (
            .in_data({
                         in_data[573],
                         in_data[722],
                         in_data[502],
                         in_data[610],
                         in_data[89],
                         in_data[192]
                    }),
            .out_data(lut_485_out)
        );

reg   lut_485_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_485_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_485_ff <= lut_485_out;
    end
end

assign out_data[485] = lut_485_ff;




// LUT : 486

wire lut_486_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110010100000001000000010010010000011110000101000000011000000),
            .DEVICE(DEVICE)
        )
    i_lut_486
        (
            .in_data({
                         in_data[101],
                         in_data[491],
                         in_data[264],
                         in_data[48],
                         in_data[612],
                         in_data[177]
                    }),
            .out_data(lut_486_out)
        );

reg   lut_486_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_486_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_486_ff <= lut_486_out;
    end
end

assign out_data[486] = lut_486_ff;




// LUT : 487

wire lut_487_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010110111101101111110110111111010100010101101101011111111110),
            .DEVICE(DEVICE)
        )
    i_lut_487
        (
            .in_data({
                         in_data[637],
                         in_data[379],
                         in_data[537],
                         in_data[660],
                         in_data[240],
                         in_data[533]
                    }),
            .out_data(lut_487_out)
        );

reg   lut_487_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_487_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_487_ff <= lut_487_out;
    end
end

assign out_data[487] = lut_487_ff;




// LUT : 488

wire lut_488_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101001011001001101010111110001011100010010110111111110000111110),
            .DEVICE(DEVICE)
        )
    i_lut_488
        (
            .in_data({
                         in_data[105],
                         in_data[617],
                         in_data[70],
                         in_data[190],
                         in_data[3],
                         in_data[754]
                    }),
            .out_data(lut_488_out)
        );

reg   lut_488_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_488_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_488_ff <= lut_488_out;
    end
end

assign out_data[488] = lut_488_ff;




// LUT : 489

wire lut_489_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101111010011100110000101110011111111110111111101111111011111),
            .DEVICE(DEVICE)
        )
    i_lut_489
        (
            .in_data({
                         in_data[538],
                         in_data[571],
                         in_data[482],
                         in_data[499],
                         in_data[39],
                         in_data[496]
                    }),
            .out_data(lut_489_out)
        );

reg   lut_489_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_489_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_489_ff <= lut_489_out;
    end
end

assign out_data[489] = lut_489_ff;




// LUT : 490

wire lut_490_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001101010110010101101111100010010110010001010011010011101101111),
            .DEVICE(DEVICE)
        )
    i_lut_490
        (
            .in_data({
                         in_data[107],
                         in_data[643],
                         in_data[49],
                         in_data[246],
                         in_data[74],
                         in_data[139]
                    }),
            .out_data(lut_490_out)
        );

reg   lut_490_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_490_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_490_ff <= lut_490_out;
    end
end

assign out_data[490] = lut_490_ff;




// LUT : 491

wire lut_491_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001111100100100011101001111111111111100001010101111111111101110),
            .DEVICE(DEVICE)
        )
    i_lut_491
        (
            .in_data({
                         in_data[299],
                         in_data[526],
                         in_data[390],
                         in_data[320],
                         in_data[270],
                         in_data[254]
                    }),
            .out_data(lut_491_out)
        );

reg   lut_491_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_491_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_491_ff <= lut_491_out;
    end
end

assign out_data[491] = lut_491_ff;




// LUT : 492

wire lut_492_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101101011000011111010111100011100101100010011101010111111000),
            .DEVICE(DEVICE)
        )
    i_lut_492
        (
            .in_data({
                         in_data[656],
                         in_data[277],
                         in_data[399],
                         in_data[550],
                         in_data[250],
                         in_data[779]
                    }),
            .out_data(lut_492_out)
        );

reg   lut_492_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_492_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_492_ff <= lut_492_out;
    end
end

assign out_data[492] = lut_492_ff;




// LUT : 493

wire lut_493_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010000101010010101010101111101000011011001010100111111011010),
            .DEVICE(DEVICE)
        )
    i_lut_493
        (
            .in_data({
                         in_data[354],
                         in_data[700],
                         in_data[670],
                         in_data[748],
                         in_data[519],
                         in_data[705]
                    }),
            .out_data(lut_493_out)
        );

reg   lut_493_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_493_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_493_ff <= lut_493_out;
    end
end

assign out_data[493] = lut_493_ff;




// LUT : 494

wire lut_494_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110000010000001010100010010101110101010101010111010001010101011),
            .DEVICE(DEVICE)
        )
    i_lut_494
        (
            .in_data({
                         in_data[719],
                         in_data[328],
                         in_data[711],
                         in_data[658],
                         in_data[630],
                         in_data[507]
                    }),
            .out_data(lut_494_out)
        );

reg   lut_494_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_494_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_494_ff <= lut_494_out;
    end
end

assign out_data[494] = lut_494_ff;




// LUT : 495

wire lut_495_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100101101010111110000100100011100011010100101101101000111000),
            .DEVICE(DEVICE)
        )
    i_lut_495
        (
            .in_data({
                         in_data[211],
                         in_data[780],
                         in_data[164],
                         in_data[300],
                         in_data[510],
                         in_data[382]
                    }),
            .out_data(lut_495_out)
        );

reg   lut_495_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_495_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_495_ff <= lut_495_out;
    end
end

assign out_data[495] = lut_495_ff;




// LUT : 496

wire lut_496_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001100110001011110110111111110011101110011110101111111101010),
            .DEVICE(DEVICE)
        )
    i_lut_496
        (
            .in_data({
                         in_data[436],
                         in_data[283],
                         in_data[487],
                         in_data[649],
                         in_data[551],
                         in_data[500]
                    }),
            .out_data(lut_496_out)
        );

reg   lut_496_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_496_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_496_ff <= lut_496_out;
    end
end

assign out_data[496] = lut_496_ff;




// LUT : 497

wire lut_497_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111100011100110010000010100010111000011110111100100000011000),
            .DEVICE(DEVICE)
        )
    i_lut_497
        (
            .in_data({
                         in_data[275],
                         in_data[24],
                         in_data[244],
                         in_data[782],
                         in_data[279],
                         in_data[161]
                    }),
            .out_data(lut_497_out)
        );

reg   lut_497_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_497_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_497_ff <= lut_497_out;
    end
end

assign out_data[497] = lut_497_ff;




// LUT : 498

wire lut_498_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111110010101000101111111011111011111111011100111010111101110),
            .DEVICE(DEVICE)
        )
    i_lut_498
        (
            .in_data({
                         in_data[286],
                         in_data[387],
                         in_data[229],
                         in_data[376],
                         in_data[677],
                         in_data[421]
                    }),
            .out_data(lut_498_out)
        );

reg   lut_498_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_498_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_498_ff <= lut_498_out;
    end
end

assign out_data[498] = lut_498_ff;




// LUT : 499

wire lut_499_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110111101000111110101111111111110101001011010100111011111110011),
            .DEVICE(DEVICE)
        )
    i_lut_499
        (
            .in_data({
                         in_data[597],
                         in_data[263],
                         in_data[232],
                         in_data[776],
                         in_data[672],
                         in_data[417]
                    }),
            .out_data(lut_499_out)
        );

reg   lut_499_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_499_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_499_ff <= lut_499_out;
    end
end

assign out_data[499] = lut_499_ff;




// LUT : 500

wire lut_500_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001111011010110001010010010100001111101001010110111100000101),
            .DEVICE(DEVICE)
        )
    i_lut_500
        (
            .in_data({
                         in_data[114],
                         in_data[432],
                         in_data[364],
                         in_data[774],
                         in_data[117],
                         in_data[337]
                    }),
            .out_data(lut_500_out)
        );

reg   lut_500_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_500_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_500_ff <= lut_500_out;
    end
end

assign out_data[500] = lut_500_ff;




// LUT : 501

wire lut_501_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011011011100110010011111100101000100101110011010010111101101),
            .DEVICE(DEVICE)
        )
    i_lut_501
        (
            .in_data({
                         in_data[202],
                         in_data[37],
                         in_data[497],
                         in_data[641],
                         in_data[141],
                         in_data[565]
                    }),
            .out_data(lut_501_out)
        );

reg   lut_501_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_501_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_501_ff <= lut_501_out;
    end
end

assign out_data[501] = lut_501_ff;




// LUT : 502

wire lut_502_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110101010001000011010110000011010011111110111101101111111111110),
            .DEVICE(DEVICE)
        )
    i_lut_502
        (
            .in_data({
                         in_data[167],
                         in_data[348],
                         in_data[683],
                         in_data[73],
                         in_data[303],
                         in_data[525]
                    }),
            .out_data(lut_502_out)
        );

reg   lut_502_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_502_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_502_ff <= lut_502_out;
    end
end

assign out_data[502] = lut_502_ff;




// LUT : 503

wire lut_503_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010110001101011100000101111111001010110111110011000111001100111),
            .DEVICE(DEVICE)
        )
    i_lut_503
        (
            .in_data({
                         in_data[265],
                         in_data[448],
                         in_data[241],
                         in_data[4],
                         in_data[490],
                         in_data[197]
                    }),
            .out_data(lut_503_out)
        );

reg   lut_503_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_503_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_503_ff <= lut_503_out;
    end
end

assign out_data[503] = lut_503_ff;




// LUT : 504

wire lut_504_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010011001110010010001111111101000010100000110101010111111010),
            .DEVICE(DEVICE)
        )
    i_lut_504
        (
            .in_data({
                         in_data[688],
                         in_data[363],
                         in_data[648],
                         in_data[235],
                         in_data[305],
                         in_data[681]
                    }),
            .out_data(lut_504_out)
        );

reg   lut_504_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_504_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_504_ff <= lut_504_out;
    end
end

assign out_data[504] = lut_504_ff;




// LUT : 505

wire lut_505_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001010001000100010000000100011001000110001011000000100000101),
            .DEVICE(DEVICE)
        )
    i_lut_505
        (
            .in_data({
                         in_data[400],
                         in_data[218],
                         in_data[266],
                         in_data[332],
                         in_data[423],
                         in_data[313]
                    }),
            .out_data(lut_505_out)
        );

reg   lut_505_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_505_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_505_ff <= lut_505_out;
    end
end

assign out_data[505] = lut_505_ff;




// LUT : 506

wire lut_506_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001110101001010011100000010100100011110110010100110101101011011),
            .DEVICE(DEVICE)
        )
    i_lut_506
        (
            .in_data({
                         in_data[90],
                         in_data[96],
                         in_data[653],
                         in_data[394],
                         in_data[579],
                         in_data[703]
                    }),
            .out_data(lut_506_out)
        );

reg   lut_506_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_506_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_506_ff <= lut_506_out;
    end
end

assign out_data[506] = lut_506_ff;




// LUT : 507

wire lut_507_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111001100001110100000110010110100101010010111000111110011011),
            .DEVICE(DEVICE)
        )
    i_lut_507
        (
            .in_data({
                         in_data[760],
                         in_data[416],
                         in_data[474],
                         in_data[168],
                         in_data[459],
                         in_data[556]
                    }),
            .out_data(lut_507_out)
        );

reg   lut_507_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_507_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_507_ff <= lut_507_out;
    end
end

assign out_data[507] = lut_507_ff;




// LUT : 508

wire lut_508_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111101101101011110110110100011101011001010100000110110110011),
            .DEVICE(DEVICE)
        )
    i_lut_508
        (
            .in_data({
                         in_data[163],
                         in_data[38],
                         in_data[30],
                         in_data[310],
                         in_data[94],
                         in_data[245]
                    }),
            .out_data(lut_508_out)
        );

reg   lut_508_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_508_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_508_ff <= lut_508_out;
    end
end

assign out_data[508] = lut_508_ff;




// LUT : 509

wire lut_509_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001111001110111100110000011000010111111111111111000100101110),
            .DEVICE(DEVICE)
        )
    i_lut_509
        (
            .in_data({
                         in_data[685],
                         in_data[430],
                         in_data[375],
                         in_data[709],
                         in_data[397],
                         in_data[370]
                    }),
            .out_data(lut_509_out)
        );

reg   lut_509_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_509_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_509_ff <= lut_509_out;
    end
end

assign out_data[509] = lut_509_ff;




// LUT : 510

wire lut_510_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111001001101011001010101111001010000101100000101001100100001),
            .DEVICE(DEVICE)
        )
    i_lut_510
        (
            .in_data({
                         in_data[505],
                         in_data[78],
                         in_data[239],
                         in_data[87],
                         in_data[158],
                         in_data[548]
                    }),
            .out_data(lut_510_out)
        );

reg   lut_510_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_510_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_510_ff <= lut_510_out;
    end
end

assign out_data[510] = lut_510_ff;




// LUT : 511

wire lut_511_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010100110101110000010001011001011110100011001000000101111100),
            .DEVICE(DEVICE)
        )
    i_lut_511
        (
            .in_data({
                         in_data[644],
                         in_data[224],
                         in_data[646],
                         in_data[479],
                         in_data[739],
                         in_data[694]
                    }),
            .out_data(lut_511_out)
        );

reg   lut_511_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_511_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_511_ff <= lut_511_out;
    end
end

assign out_data[511] = lut_511_ff;




// LUT : 512

wire lut_512_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111110100010011000100010001110011001110110001010111011101),
            .DEVICE(DEVICE)
        )
    i_lut_512
        (
            .in_data({
                         in_data[159],
                         in_data[710],
                         in_data[380],
                         in_data[625],
                         in_data[20],
                         in_data[636]
                    }),
            .out_data(lut_512_out)
        );

reg   lut_512_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_512_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_512_ff <= lut_512_out;
    end
end

assign out_data[512] = lut_512_ff;




// LUT : 513

wire lut_513_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001111000101001000011010000000010111100001101011100111111100011),
            .DEVICE(DEVICE)
        )
    i_lut_513
        (
            .in_data({
                         in_data[166],
                         in_data[667],
                         in_data[408],
                         in_data[607],
                         in_data[195],
                         in_data[541]
                    }),
            .out_data(lut_513_out)
        );

reg   lut_513_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_513_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_513_ff <= lut_513_out;
    end
end

assign out_data[513] = lut_513_ff;




// LUT : 514

wire lut_514_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111010000111101111111101111110111000100101000010011100110000),
            .DEVICE(DEVICE)
        )
    i_lut_514
        (
            .in_data({
                         in_data[52],
                         in_data[708],
                         in_data[572],
                         in_data[88],
                         in_data[296],
                         in_data[713]
                    }),
            .out_data(lut_514_out)
        );

reg   lut_514_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_514_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_514_ff <= lut_514_out;
    end
end

assign out_data[514] = lut_514_ff;




// LUT : 515

wire lut_515_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111010000000011101110110011100101100011001000000010111111101),
            .DEVICE(DEVICE)
        )
    i_lut_515
        (
            .in_data({
                         in_data[598],
                         in_data[71],
                         in_data[186],
                         in_data[698],
                         in_data[373],
                         in_data[412]
                    }),
            .out_data(lut_515_out)
        );

reg   lut_515_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_515_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_515_ff <= lut_515_out;
    end
end

assign out_data[515] = lut_515_ff;




// LUT : 516

wire lut_516_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001110110100011111101000101000011110111001100010010101001000010),
            .DEVICE(DEVICE)
        )
    i_lut_516
        (
            .in_data({
                         in_data[772],
                         in_data[61],
                         in_data[324],
                         in_data[31],
                         in_data[200],
                         in_data[451]
                    }),
            .out_data(lut_516_out)
        );

reg   lut_516_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_516_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_516_ff <= lut_516_out;
    end
end

assign out_data[516] = lut_516_ff;




// LUT : 517

wire lut_517_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100010111011101000010110010111001111100011110001101010011010),
            .DEVICE(DEVICE)
        )
    i_lut_517
        (
            .in_data({
                         in_data[769],
                         in_data[230],
                         in_data[152],
                         in_data[9],
                         in_data[404],
                         in_data[149]
                    }),
            .out_data(lut_517_out)
        );

reg   lut_517_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_517_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_517_ff <= lut_517_out;
    end
end

assign out_data[517] = lut_517_ff;




// LUT : 518

wire lut_518_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010110011101000011000101111111110011000110000011100001011111111),
            .DEVICE(DEVICE)
        )
    i_lut_518
        (
            .in_data({
                         in_data[524],
                         in_data[485],
                         in_data[85],
                         in_data[469],
                         in_data[106],
                         in_data[123]
                    }),
            .out_data(lut_518_out)
        );

reg   lut_518_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_518_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_518_ff <= lut_518_out;
    end
end

assign out_data[518] = lut_518_ff;




// LUT : 519

wire lut_519_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001011101111100000000010100001010011111010001001100011111011000),
            .DEVICE(DEVICE)
        )
    i_lut_519
        (
            .in_data({
                         in_data[456],
                         in_data[243],
                         in_data[621],
                         in_data[18],
                         in_data[109],
                         in_data[84]
                    }),
            .out_data(lut_519_out)
        );

reg   lut_519_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_519_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_519_ff <= lut_519_out;
    end
end

assign out_data[519] = lut_519_ff;




// LUT : 520

wire lut_520_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100010100010010000111000000000000100110111000100001101010011),
            .DEVICE(DEVICE)
        )
    i_lut_520
        (
            .in_data({
                         in_data[401],
                         in_data[51],
                         in_data[153],
                         in_data[559],
                         in_data[473],
                         in_data[600]
                    }),
            .out_data(lut_520_out)
        );

reg   lut_520_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_520_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_520_ff <= lut_520_out;
    end
end

assign out_data[520] = lut_520_ff;




// LUT : 521

wire lut_521_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110000000100110010010101100110110000101011001111011000011111111),
            .DEVICE(DEVICE)
        )
    i_lut_521
        (
            .in_data({
                         in_data[279],
                         in_data[703],
                         in_data[777],
                         in_data[733],
                         in_data[561],
                         in_data[53]
                    }),
            .out_data(lut_521_out)
        );

reg   lut_521_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_521_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_521_ff <= lut_521_out;
    end
end

assign out_data[521] = lut_521_ff;




// LUT : 522

wire lut_522_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010101010101110010111011011110101011011100011111001001110010),
            .DEVICE(DEVICE)
        )
    i_lut_522
        (
            .in_data({
                         in_data[358],
                         in_data[504],
                         in_data[13],
                         in_data[474],
                         in_data[385],
                         in_data[641]
                    }),
            .out_data(lut_522_out)
        );

reg   lut_522_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_522_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_522_ff <= lut_522_out;
    end
end

assign out_data[522] = lut_522_ff;




// LUT : 523

wire lut_523_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110110111111011111010010110100100001100000010011000101001101),
            .DEVICE(DEVICE)
        )
    i_lut_523
        (
            .in_data({
                         in_data[497],
                         in_data[573],
                         in_data[314],
                         in_data[306],
                         in_data[454],
                         in_data[405]
                    }),
            .out_data(lut_523_out)
        );

reg   lut_523_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_523_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_523_ff <= lut_523_out;
    end
end

assign out_data[523] = lut_523_ff;




// LUT : 524

wire lut_524_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011011001000001101101010000001000000000000001100011001001001),
            .DEVICE(DEVICE)
        )
    i_lut_524
        (
            .in_data({
                         in_data[669],
                         in_data[155],
                         in_data[14],
                         in_data[148],
                         in_data[770],
                         in_data[557]
                    }),
            .out_data(lut_524_out)
        );

reg   lut_524_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_524_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_524_ff <= lut_524_out;
    end
end

assign out_data[524] = lut_524_ff;




// LUT : 525

wire lut_525_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011011110101111101111011101111100000010100011111011100111110),
            .DEVICE(DEVICE)
        )
    i_lut_525
        (
            .in_data({
                         in_data[161],
                         in_data[138],
                         in_data[686],
                         in_data[667],
                         in_data[21],
                         in_data[460]
                    }),
            .out_data(lut_525_out)
        );

reg   lut_525_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_525_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_525_ff <= lut_525_out;
    end
end

assign out_data[525] = lut_525_ff;




// LUT : 526

wire lut_526_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111110101111011111110011111111111111111111110000101011111111),
            .DEVICE(DEVICE)
        )
    i_lut_526
        (
            .in_data({
                         in_data[67],
                         in_data[243],
                         in_data[490],
                         in_data[247],
                         in_data[376],
                         in_data[550]
                    }),
            .out_data(lut_526_out)
        );

reg   lut_526_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_526_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_526_ff <= lut_526_out;
    end
end

assign out_data[526] = lut_526_ff;




// LUT : 527

wire lut_527_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010000011011010100110110000001100111000111100011101101101110),
            .DEVICE(DEVICE)
        )
    i_lut_527
        (
            .in_data({
                         in_data[17],
                         in_data[710],
                         in_data[638],
                         in_data[606],
                         in_data[419],
                         in_data[107]
                    }),
            .out_data(lut_527_out)
        );

reg   lut_527_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_527_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_527_ff <= lut_527_out;
    end
end

assign out_data[527] = lut_527_ff;




// LUT : 528

wire lut_528_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101001110111011101000000000010110110110101111111001100000001111),
            .DEVICE(DEVICE)
        )
    i_lut_528
        (
            .in_data({
                         in_data[574],
                         in_data[700],
                         in_data[422],
                         in_data[99],
                         in_data[514],
                         in_data[555]
                    }),
            .out_data(lut_528_out)
        );

reg   lut_528_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_528_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_528_ff <= lut_528_out;
    end
end

assign out_data[528] = lut_528_ff;




// LUT : 529

wire lut_529_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111101010100011111111000010011000010101111000100101100011101),
            .DEVICE(DEVICE)
        )
    i_lut_529
        (
            .in_data({
                         in_data[298],
                         in_data[109],
                         in_data[529],
                         in_data[713],
                         in_data[23],
                         in_data[255]
                    }),
            .out_data(lut_529_out)
        );

reg   lut_529_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_529_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_529_ff <= lut_529_out;
    end
end

assign out_data[529] = lut_529_ff;




// LUT : 530

wire lut_530_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000110100000011111100000111100000001110001110001100111100100000),
            .DEVICE(DEVICE)
        )
    i_lut_530
        (
            .in_data({
                         in_data[285],
                         in_data[640],
                         in_data[636],
                         in_data[44],
                         in_data[120],
                         in_data[477]
                    }),
            .out_data(lut_530_out)
        );

reg   lut_530_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_530_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_530_ff <= lut_530_out;
    end
end

assign out_data[530] = lut_530_ff;




// LUT : 531

wire lut_531_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001010000000011010111010010010000001011011100100110010110011),
            .DEVICE(DEVICE)
        )
    i_lut_531
        (
            .in_data({
                         in_data[509],
                         in_data[633],
                         in_data[614],
                         in_data[412],
                         in_data[7],
                         in_data[396]
                    }),
            .out_data(lut_531_out)
        );

reg   lut_531_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_531_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_531_ff <= lut_531_out;
    end
end

assign out_data[531] = lut_531_ff;




// LUT : 532

wire lut_532_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100111111101110111000111111011100101110001011001110001010100),
            .DEVICE(DEVICE)
        )
    i_lut_532
        (
            .in_data({
                         in_data[235],
                         in_data[513],
                         in_data[371],
                         in_data[167],
                         in_data[558],
                         in_data[4]
                    }),
            .out_data(lut_532_out)
        );

reg   lut_532_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_532_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_532_ff <= lut_532_out;
    end
end

assign out_data[532] = lut_532_ff;




// LUT : 533

wire lut_533_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011110101111001011111000111101010111111000111110011111010010),
            .DEVICE(DEVICE)
        )
    i_lut_533
        (
            .in_data({
                         in_data[172],
                         in_data[597],
                         in_data[173],
                         in_data[45],
                         in_data[714],
                         in_data[119]
                    }),
            .out_data(lut_533_out)
        );

reg   lut_533_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_533_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_533_ff <= lut_533_out;
    end
end

assign out_data[533] = lut_533_ff;




// LUT : 534

wire lut_534_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010111000111000000100000010110011101110100000011111101011010),
            .DEVICE(DEVICE)
        )
    i_lut_534
        (
            .in_data({
                         in_data[5],
                         in_data[206],
                         in_data[404],
                         in_data[3],
                         in_data[301],
                         in_data[217]
                    }),
            .out_data(lut_534_out)
        );

reg   lut_534_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_534_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_534_ff <= lut_534_out;
    end
end

assign out_data[534] = lut_534_ff;




// LUT : 535

wire lut_535_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010001011010010010001010100100110010010101000110010110000001),
            .DEVICE(DEVICE)
        )
    i_lut_535
        (
            .in_data({
                         in_data[244],
                         in_data[593],
                         in_data[635],
                         in_data[169],
                         in_data[673],
                         in_data[725]
                    }),
            .out_data(lut_535_out)
        );

reg   lut_535_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_535_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_535_ff <= lut_535_out;
    end
end

assign out_data[535] = lut_535_ff;




// LUT : 536

wire lut_536_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111101111100101000010010000111011011001110001111101101111011),
            .DEVICE(DEVICE)
        )
    i_lut_536
        (
            .in_data({
                         in_data[761],
                         in_data[718],
                         in_data[519],
                         in_data[771],
                         in_data[688],
                         in_data[194]
                    }),
            .out_data(lut_536_out)
        );

reg   lut_536_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_536_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_536_ff <= lut_536_out;
    end
end

assign out_data[536] = lut_536_ff;




// LUT : 537

wire lut_537_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100110010000110010100000111111010111101111110101111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_537
        (
            .in_data({
                         in_data[253],
                         in_data[393],
                         in_data[333],
                         in_data[530],
                         in_data[494],
                         in_data[342]
                    }),
            .out_data(lut_537_out)
        );

reg   lut_537_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_537_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_537_ff <= lut_537_out;
    end
end

assign out_data[537] = lut_537_ff;




// LUT : 538

wire lut_538_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111100011110000011101001111001110101111111010000001010111100011),
            .DEVICE(DEVICE)
        )
    i_lut_538
        (
            .in_data({
                         in_data[551],
                         in_data[466],
                         in_data[390],
                         in_data[351],
                         in_data[227],
                         in_data[540]
                    }),
            .out_data(lut_538_out)
        );

reg   lut_538_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_538_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_538_ff <= lut_538_out;
    end
end

assign out_data[538] = lut_538_ff;




// LUT : 539

wire lut_539_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110011011100010100100010111100111111011111111011001101011101),
            .DEVICE(DEVICE)
        )
    i_lut_539
        (
            .in_data({
                         in_data[541],
                         in_data[426],
                         in_data[757],
                         in_data[632],
                         in_data[705],
                         in_data[31]
                    }),
            .out_data(lut_539_out)
        );

reg   lut_539_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_539_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_539_ff <= lut_539_out;
    end
end

assign out_data[539] = lut_539_ff;




// LUT : 540

wire lut_540_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111110100011010110011100000110001010000100011000111001100111),
            .DEVICE(DEVICE)
        )
    i_lut_540
        (
            .in_data({
                         in_data[40],
                         in_data[444],
                         in_data[736],
                         in_data[470],
                         in_data[642],
                         in_data[162]
                    }),
            .out_data(lut_540_out)
        );

reg   lut_540_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_540_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_540_ff <= lut_540_out;
    end
end

assign out_data[540] = lut_540_ff;




// LUT : 541

wire lut_541_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010001111111101000000011000010100101101011111010011110101110),
            .DEVICE(DEVICE)
        )
    i_lut_541
        (
            .in_data({
                         in_data[453],
                         in_data[408],
                         in_data[296],
                         in_data[395],
                         in_data[457],
                         in_data[359]
                    }),
            .out_data(lut_541_out)
        );

reg   lut_541_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_541_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_541_ff <= lut_541_out;
    end
end

assign out_data[541] = lut_541_ff;




// LUT : 542

wire lut_542_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110010111110110100110001000111100100100001111101010111111010),
            .DEVICE(DEVICE)
        )
    i_lut_542
        (
            .in_data({
                         in_data[15],
                         in_data[349],
                         in_data[488],
                         in_data[37],
                         in_data[543],
                         in_data[379]
                    }),
            .out_data(lut_542_out)
        );

reg   lut_542_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_542_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_542_ff <= lut_542_out;
    end
end

assign out_data[542] = lut_542_ff;




// LUT : 543

wire lut_543_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000110111000001101010110010100011111011000100101000101010101),
            .DEVICE(DEVICE)
        )
    i_lut_543
        (
            .in_data({
                         in_data[199],
                         in_data[448],
                         in_data[462],
                         in_data[368],
                         in_data[441],
                         in_data[327]
                    }),
            .out_data(lut_543_out)
        );

reg   lut_543_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_543_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_543_ff <= lut_543_out;
    end
end

assign out_data[543] = lut_543_ff;




// LUT : 544

wire lut_544_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010100100001101110001011111000101010010010011000001111111100),
            .DEVICE(DEVICE)
        )
    i_lut_544
        (
            .in_data({
                         in_data[249],
                         in_data[281],
                         in_data[752],
                         in_data[521],
                         in_data[527],
                         in_data[322]
                    }),
            .out_data(lut_544_out)
        );

reg   lut_544_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_544_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_544_ff <= lut_544_out;
    end
end

assign out_data[544] = lut_544_ff;




// LUT : 545

wire lut_545_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100011011010110111011010010101010010000110000110110100000101),
            .DEVICE(DEVICE)
        )
    i_lut_545
        (
            .in_data({
                         in_data[476],
                         in_data[12],
                         in_data[589],
                         in_data[370],
                         in_data[213],
                         in_data[94]
                    }),
            .out_data(lut_545_out)
        );

reg   lut_545_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_545_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_545_ff <= lut_545_out;
    end
end

assign out_data[545] = lut_545_ff;




// LUT : 546

wire lut_546_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111100000001101001011001000110100001000011001000100110011111101),
            .DEVICE(DEVICE)
        )
    i_lut_546
        (
            .in_data({
                         in_data[299],
                         in_data[373],
                         in_data[38],
                         in_data[49],
                         in_data[242],
                         in_data[417]
                    }),
            .out_data(lut_546_out)
        );

reg   lut_546_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_546_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_546_ff <= lut_546_out;
    end
end

assign out_data[546] = lut_546_ff;




// LUT : 547

wire lut_547_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000111000100100001010001100111111110011000010111100100101011),
            .DEVICE(DEVICE)
        )
    i_lut_547
        (
            .in_data({
                         in_data[318],
                         in_data[225],
                         in_data[450],
                         in_data[2],
                         in_data[278],
                         in_data[414]
                    }),
            .out_data(lut_547_out)
        );

reg   lut_547_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_547_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_547_ff <= lut_547_out;
    end
end

assign out_data[547] = lut_547_ff;




// LUT : 548

wire lut_548_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001111011010110110001000101010001101001001001111010110101100),
            .DEVICE(DEVICE)
        )
    i_lut_548
        (
            .in_data({
                         in_data[696],
                         in_data[582],
                         in_data[357],
                         in_data[277],
                         in_data[292],
                         in_data[780]
                    }),
            .out_data(lut_548_out)
        );

reg   lut_548_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_548_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_548_ff <= lut_548_out;
    end
end

assign out_data[548] = lut_548_ff;




// LUT : 549

wire lut_549_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000110000111001110010101111111110111001011111111010000100010),
            .DEVICE(DEVICE)
        )
    i_lut_549
        (
            .in_data({
                         in_data[617],
                         in_data[241],
                         in_data[493],
                         in_data[240],
                         in_data[92],
                         in_data[297]
                    }),
            .out_data(lut_549_out)
        );

reg   lut_549_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_549_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_549_ff <= lut_549_out;
    end
end

assign out_data[549] = lut_549_ff;




// LUT : 550

wire lut_550_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010010010000101000001101110011110000001101011000000001010111),
            .DEVICE(DEVICE)
        )
    i_lut_550
        (
            .in_data({
                         in_data[501],
                         in_data[384],
                         in_data[147],
                         in_data[479],
                         in_data[622],
                         in_data[528]
                    }),
            .out_data(lut_550_out)
        );

reg   lut_550_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_550_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_550_ff <= lut_550_out;
    end
end

assign out_data[550] = lut_550_ff;




// LUT : 551

wire lut_551_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011110101111111101011110111010111101101010101011111110111110),
            .DEVICE(DEVICE)
        )
    i_lut_551
        (
            .in_data({
                         in_data[160],
                         in_data[525],
                         in_data[435],
                         in_data[680],
                         in_data[689],
                         in_data[704]
                    }),
            .out_data(lut_551_out)
        );

reg   lut_551_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_551_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_551_ff <= lut_551_out;
    end
end

assign out_data[551] = lut_551_ff;




// LUT : 552

wire lut_552_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000100000100011100000011001101111111100000000100110000000011),
            .DEVICE(DEVICE)
        )
    i_lut_552
        (
            .in_data({
                         in_data[246],
                         in_data[133],
                         in_data[674],
                         in_data[332],
                         in_data[250],
                         in_data[291]
                    }),
            .out_data(lut_552_out)
        );

reg   lut_552_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_552_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_552_ff <= lut_552_out;
    end
end

assign out_data[552] = lut_552_ff;




// LUT : 553

wire lut_553_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010111101001111110001111001110000101011100001111110011110011101),
            .DEVICE(DEVICE)
        )
    i_lut_553
        (
            .in_data({
                         in_data[730],
                         in_data[142],
                         in_data[562],
                         in_data[694],
                         in_data[679],
                         in_data[273]
                    }),
            .out_data(lut_553_out)
        );

reg   lut_553_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_553_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_553_ff <= lut_553_out;
    end
end

assign out_data[553] = lut_553_ff;




// LUT : 554

wire lut_554_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111100110010010001100111100110011010001100100001110011101011111),
            .DEVICE(DEVICE)
        )
    i_lut_554
        (
            .in_data({
                         in_data[566],
                         in_data[707],
                         in_data[168],
                         in_data[309],
                         in_data[533],
                         in_data[445]
                    }),
            .out_data(lut_554_out)
        );

reg   lut_554_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_554_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_554_ff <= lut_554_out;
    end
end

assign out_data[554] = lut_554_ff;




// LUT : 555

wire lut_555_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001010110111111011001111100010100101111110010011111101001010),
            .DEVICE(DEVICE)
        )
    i_lut_555
        (
            .in_data({
                         in_data[701],
                         in_data[166],
                         in_data[744],
                         in_data[664],
                         in_data[418],
                         in_data[340]
                    }),
            .out_data(lut_555_out)
        );

reg   lut_555_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_555_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_555_ff <= lut_555_out;
    end
end

assign out_data[555] = lut_555_ff;




// LUT : 556

wire lut_556_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001011000000001000110100001101001111011010010110010101000011),
            .DEVICE(DEVICE)
        )
    i_lut_556
        (
            .in_data({
                         in_data[186],
                         in_data[130],
                         in_data[719],
                         in_data[536],
                         in_data[65],
                         in_data[495]
                    }),
            .out_data(lut_556_out)
        );

reg   lut_556_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_556_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_556_ff <= lut_556_out;
    end
end

assign out_data[556] = lut_556_ff;




// LUT : 557

wire lut_557_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110101101111111011011101000010111011100001010000000010001100),
            .DEVICE(DEVICE)
        )
    i_lut_557
        (
            .in_data({
                         in_data[724],
                         in_data[85],
                         in_data[135],
                         in_data[60],
                         in_data[583],
                         in_data[100]
                    }),
            .out_data(lut_557_out)
        );

reg   lut_557_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_557_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_557_ff <= lut_557_out;
    end
end

assign out_data[557] = lut_557_ff;




// LUT : 558

wire lut_558_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101010011001011111111111111110000110110010110101001111111111),
            .DEVICE(DEVICE)
        )
    i_lut_558
        (
            .in_data({
                         in_data[402],
                         in_data[54],
                         in_data[268],
                         in_data[128],
                         in_data[378],
                         in_data[212]
                    }),
            .out_data(lut_558_out)
        );

reg   lut_558_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_558_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_558_ff <= lut_558_out;
    end
end

assign out_data[558] = lut_558_ff;




// LUT : 559

wire lut_559_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001011111111101111101111111100110000110010100100011111000111),
            .DEVICE(DEVICE)
        )
    i_lut_559
        (
            .in_data({
                         in_data[443],
                         in_data[690],
                         in_data[538],
                         in_data[579],
                         in_data[41],
                         in_data[482]
                    }),
            .out_data(lut_559_out)
        );

reg   lut_559_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_559_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_559_ff <= lut_559_out;
    end
end

assign out_data[559] = lut_559_ff;




// LUT : 560

wire lut_560_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110110000110010000110010001101011011100000001001110100000110100),
            .DEVICE(DEVICE)
        )
    i_lut_560
        (
            .in_data({
                         in_data[723],
                         in_data[548],
                         in_data[364],
                         in_data[756],
                         in_data[429],
                         in_data[123]
                    }),
            .out_data(lut_560_out)
        );

reg   lut_560_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_560_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_560_ff <= lut_560_out;
    end
end

assign out_data[560] = lut_560_ff;




// LUT : 561

wire lut_561_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011011001111101111011001111010011010111011101000101110111111000),
            .DEVICE(DEVICE)
        )
    i_lut_561
        (
            .in_data({
                         in_data[215],
                         in_data[415],
                         in_data[70],
                         in_data[542],
                         in_data[136],
                         in_data[678]
                    }),
            .out_data(lut_561_out)
        );

reg   lut_561_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_561_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_561_ff <= lut_561_out;
    end
end

assign out_data[561] = lut_561_ff;




// LUT : 562

wire lut_562_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001100100111001000001010010000011111011011000000001001001000100),
            .DEVICE(DEVICE)
        )
    i_lut_562
        (
            .in_data({
                         in_data[449],
                         in_data[745],
                         in_data[760],
                         in_data[308],
                         in_data[407],
                         in_data[776]
                    }),
            .out_data(lut_562_out)
        );

reg   lut_562_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_562_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_562_ff <= lut_562_out;
    end
end

assign out_data[562] = lut_562_ff;




// LUT : 563

wire lut_563_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000001110100011000011010100000010010000000110100001100000011),
            .DEVICE(DEVICE)
        )
    i_lut_563
        (
            .in_data({
                         in_data[734],
                         in_data[461],
                         in_data[360],
                         in_data[423],
                         in_data[621],
                         in_data[329]
                    }),
            .out_data(lut_563_out)
        );

reg   lut_563_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_563_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_563_ff <= lut_563_out;
    end
end

assign out_data[563] = lut_563_ff;




// LUT : 564

wire lut_564_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000000001000010000110100110000000110000000000000000001011100),
            .DEVICE(DEVICE)
        )
    i_lut_564
        (
            .in_data({
                         in_data[498],
                         in_data[122],
                         in_data[506],
                         in_data[569],
                         in_data[567],
                         in_data[455]
                    }),
            .out_data(lut_564_out)
        );

reg   lut_564_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_564_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_564_ff <= lut_564_out;
    end
end

assign out_data[564] = lut_564_ff;




// LUT : 565

wire lut_565_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000001000110001101101011100001010100001001011000110000011010),
            .DEVICE(DEVICE)
        )
    i_lut_565
        (
            .in_data({
                         in_data[425],
                         in_data[502],
                         in_data[708],
                         in_data[63],
                         in_data[372],
                         in_data[197]
                    }),
            .out_data(lut_565_out)
        );

reg   lut_565_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_565_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_565_ff <= lut_565_out;
    end
end

assign out_data[565] = lut_565_ff;




// LUT : 566

wire lut_566_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001100010101101101110101100001100000000101110101101100101111111),
            .DEVICE(DEVICE)
        )
    i_lut_566
        (
            .in_data({
                         in_data[59],
                         in_data[205],
                         in_data[468],
                         in_data[531],
                         in_data[742],
                         in_data[272]
                    }),
            .out_data(lut_566_out)
        );

reg   lut_566_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_566_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_566_ff <= lut_566_out;
    end
end

assign out_data[566] = lut_566_ff;




// LUT : 567

wire lut_567_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001110001011010100010000001000011010001011111010100001000010110),
            .DEVICE(DEVICE)
        )
    i_lut_567
        (
            .in_data({
                         in_data[264],
                         in_data[88],
                         in_data[183],
                         in_data[524],
                         in_data[388],
                         in_data[492]
                    }),
            .out_data(lut_567_out)
        );

reg   lut_567_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_567_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_567_ff <= lut_567_out;
    end
end

assign out_data[567] = lut_567_ff;




// LUT : 568

wire lut_568_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100101111111111010101001010100000000000000110101110101110101),
            .DEVICE(DEVICE)
        )
    i_lut_568
        (
            .in_data({
                         in_data[112],
                         in_data[76],
                         in_data[438],
                         in_data[601],
                         in_data[157],
                         in_data[439]
                    }),
            .out_data(lut_568_out)
        );

reg   lut_568_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_568_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_568_ff <= lut_568_out;
    end
end

assign out_data[568] = lut_568_ff;




// LUT : 569

wire lut_569_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110111011101101110101011101110010100110111011011110111111111),
            .DEVICE(DEVICE)
        )
    i_lut_569
        (
            .in_data({
                         in_data[326],
                         in_data[229],
                         in_data[749],
                         in_data[545],
                         in_data[339],
                         in_data[259]
                    }),
            .out_data(lut_569_out)
        );

reg   lut_569_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_569_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_569_ff <= lut_569_out;
    end
end

assign out_data[569] = lut_569_ff;




// LUT : 570

wire lut_570_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010011000100001000011110100001010111001100110100110111110100110),
            .DEVICE(DEVICE)
        )
    i_lut_570
        (
            .in_data({
                         in_data[9],
                         in_data[68],
                         in_data[374],
                         in_data[475],
                         in_data[113],
                         in_data[275]
                    }),
            .out_data(lut_570_out)
        );

reg   lut_570_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_570_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_570_ff <= lut_570_out;
    end
end

assign out_data[570] = lut_570_ff;




// LUT : 571

wire lut_571_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000011100000010001001010100000100000010010110111110001111111),
            .DEVICE(DEVICE)
        )
    i_lut_571
        (
            .in_data({
                         in_data[300],
                         in_data[591],
                         in_data[544],
                         in_data[767],
                         in_data[687],
                         in_data[434]
                    }),
            .out_data(lut_571_out)
        );

reg   lut_571_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_571_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_571_ff <= lut_571_out;
    end
end

assign out_data[571] = lut_571_ff;




// LUT : 572

wire lut_572_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001001110000110011111100110000001011101101110110011111010110010),
            .DEVICE(DEVICE)
        )
    i_lut_572
        (
            .in_data({
                         in_data[537],
                         in_data[549],
                         in_data[615],
                         in_data[338],
                         in_data[295],
                         in_data[684]
                    }),
            .out_data(lut_572_out)
        );

reg   lut_572_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_572_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_572_ff <= lut_572_out;
    end
end

assign out_data[572] = lut_572_ff;




// LUT : 573

wire lut_573_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000100110001000100000001000101110101001110000100101100011001),
            .DEVICE(DEVICE)
        )
    i_lut_573
        (
            .in_data({
                         in_data[575],
                         in_data[198],
                         in_data[584],
                         in_data[383],
                         in_data[552],
                         in_data[702]
                    }),
            .out_data(lut_573_out)
        );

reg   lut_573_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_573_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_573_ff <= lut_573_out;
    end
end

assign out_data[573] = lut_573_ff;




// LUT : 574

wire lut_574_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001011010100010110111010100010000001110010010110111110101110111),
            .DEVICE(DEVICE)
        )
    i_lut_574
        (
            .in_data({
                         in_data[293],
                         in_data[84],
                         in_data[177],
                         in_data[483],
                         in_data[263],
                         in_data[345]
                    }),
            .out_data(lut_574_out)
        );

reg   lut_574_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_574_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_574_ff <= lut_574_out;
    end
end

assign out_data[574] = lut_574_ff;




// LUT : 575

wire lut_575_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000111010110101110101010011111011101111001101100010011001100),
            .DEVICE(DEVICE)
        )
    i_lut_575
        (
            .in_data({
                         in_data[252],
                         in_data[18],
                         in_data[467],
                         in_data[739],
                         in_data[324],
                         in_data[740]
                    }),
            .out_data(lut_575_out)
        );

reg   lut_575_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_575_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_575_ff <= lut_575_out;
    end
end

assign out_data[575] = lut_575_ff;




// LUT : 576

wire lut_576_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001111110011010110001111001100111101001111000101001101110111),
            .DEVICE(DEVICE)
        )
    i_lut_576
        (
            .in_data({
                         in_data[489],
                         in_data[754],
                         in_data[728],
                         in_data[682],
                         in_data[697],
                         in_data[81]
                    }),
            .out_data(lut_576_out)
        );

reg   lut_576_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_576_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_576_ff <= lut_576_out;
    end
end

assign out_data[576] = lut_576_ff;




// LUT : 577

wire lut_577_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001100110011101110001000100010110111101111111111011100101000),
            .DEVICE(DEVICE)
        )
    i_lut_577
        (
            .in_data({
                         in_data[353],
                         in_data[102],
                         in_data[218],
                         in_data[628],
                         in_data[392],
                         in_data[623]
                    }),
            .out_data(lut_577_out)
        );

reg   lut_577_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_577_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_577_ff <= lut_577_out;
    end
end

assign out_data[577] = lut_577_ff;




// LUT : 578

wire lut_578_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000100101101010101110100110001111010010100101000101010100000),
            .DEVICE(DEVICE)
        )
    i_lut_578
        (
            .in_data({
                         in_data[311],
                         in_data[22],
                         in_data[608],
                         in_data[656],
                         in_data[485],
                         in_data[305]
                    }),
            .out_data(lut_578_out)
        );

reg   lut_578_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_578_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_578_ff <= lut_578_out;
    end
end

assign out_data[578] = lut_578_ff;




// LUT : 579

wire lut_579_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010111100001010110110000000010100011000101001001101110110000),
            .DEVICE(DEVICE)
        )
    i_lut_579
        (
            .in_data({
                         in_data[465],
                         in_data[224],
                         in_data[346],
                         in_data[699],
                         in_data[95],
                         in_data[207]
                    }),
            .out_data(lut_579_out)
        );

reg   lut_579_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_579_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_579_ff <= lut_579_out;
    end
end

assign out_data[579] = lut_579_ff;




// LUT : 580

wire lut_580_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001101101000100110001000100010001001111010001001111101000000101),
            .DEVICE(DEVICE)
        )
    i_lut_580
        (
            .in_data({
                         in_data[625],
                         in_data[565],
                         in_data[334],
                         in_data[440],
                         in_data[380],
                         in_data[96]
                    }),
            .out_data(lut_580_out)
        );

reg   lut_580_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_580_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_580_ff <= lut_580_out;
    end
end

assign out_data[580] = lut_580_ff;




// LUT : 581

wire lut_581_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110101001111111110001001101111110100001110111111110101011101110),
            .DEVICE(DEVICE)
        )
    i_lut_581
        (
            .in_data({
                         in_data[151],
                         in_data[580],
                         in_data[27],
                         in_data[683],
                         in_data[262],
                         in_data[121]
                    }),
            .out_data(lut_581_out)
        );

reg   lut_581_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_581_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_581_ff <= lut_581_out;
    end
end

assign out_data[581] = lut_581_ff;




// LUT : 582

wire lut_582_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001001000111000011001000011111011011001100010001101111011100),
            .DEVICE(DEVICE)
        )
    i_lut_582
        (
            .in_data({
                         in_data[643],
                         in_data[768],
                         in_data[775],
                         in_data[261],
                         in_data[646],
                         in_data[594]
                    }),
            .out_data(lut_582_out)
        );

reg   lut_582_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_582_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_582_ff <= lut_582_out;
    end
end

assign out_data[582] = lut_582_ff;




// LUT : 583

wire lut_583_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001100000000010100000010111000010111100110110000001000001110011),
            .DEVICE(DEVICE)
        )
    i_lut_583
        (
            .in_data({
                         in_data[751],
                         in_data[491],
                         in_data[79],
                         in_data[534],
                         in_data[698],
                         in_data[663]
                    }),
            .out_data(lut_583_out)
        );

reg   lut_583_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_583_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_583_ff <= lut_583_out;
    end
end

assign out_data[583] = lut_583_ff;




// LUT : 584

wire lut_584_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001100100110001100011010011110001101011111111001100111100111100),
            .DEVICE(DEVICE)
        )
    i_lut_584
        (
            .in_data({
                         in_data[269],
                         in_data[657],
                         in_data[39],
                         in_data[766],
                         in_data[114],
                         in_data[712]
                    }),
            .out_data(lut_584_out)
        );

reg   lut_584_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_584_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_584_ff <= lut_584_out;
    end
end

assign out_data[584] = lut_584_ff;




// LUT : 585

wire lut_585_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010100101101100010000010111000101101001010001000100001010101),
            .DEVICE(DEVICE)
        )
    i_lut_585
        (
            .in_data({
                         in_data[189],
                         in_data[753],
                         in_data[499],
                         in_data[209],
                         in_data[381],
                         in_data[362]
                    }),
            .out_data(lut_585_out)
        );

reg   lut_585_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_585_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_585_ff <= lut_585_out;
    end
end

assign out_data[585] = lut_585_ff;




// LUT : 586

wire lut_586_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001100101111010000011111000101010010111100001100110011110000),
            .DEVICE(DEVICE)
        )
    i_lut_586
        (
            .in_data({
                         in_data[350],
                         in_data[176],
                         in_data[336],
                         in_data[738],
                         in_data[331],
                         in_data[458]
                    }),
            .out_data(lut_586_out)
        );

reg   lut_586_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_586_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_586_ff <= lut_586_out;
    end
end

assign out_data[586] = lut_586_ff;




// LUT : 587

wire lut_587_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001110100010111001010000000001111000101000101011110000110011),
            .DEVICE(DEVICE)
        )
    i_lut_587
        (
            .in_data({
                         in_data[188],
                         in_data[321],
                         in_data[764],
                         in_data[203],
                         in_data[639],
                         in_data[546]
                    }),
            .out_data(lut_587_out)
        );

reg   lut_587_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_587_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_587_ff <= lut_587_out;
    end
end

assign out_data[587] = lut_587_ff;




// LUT : 588

wire lut_588_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000001110001111110011011001011000100001001111001010110110011),
            .DEVICE(DEVICE)
        )
    i_lut_588
        (
            .in_data({
                         in_data[662],
                         in_data[146],
                         in_data[62],
                         in_data[317],
                         in_data[722],
                         in_data[230]
                    }),
            .out_data(lut_588_out)
        );

reg   lut_588_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_588_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_588_ff <= lut_588_out;
    end
end

assign out_data[588] = lut_588_ff;




// LUT : 589

wire lut_589_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011010001001001000011100111100100110100010011000011111111110111),
            .DEVICE(DEVICE)
        )
    i_lut_589
        (
            .in_data({
                         in_data[741],
                         in_data[563],
                         in_data[73],
                         in_data[400],
                         in_data[46],
                         in_data[50]
                    }),
            .out_data(lut_589_out)
        );

reg   lut_589_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_589_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_589_ff <= lut_589_out;
    end
end

assign out_data[589] = lut_589_ff;




// LUT : 590

wire lut_590_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100001101000000101111100001101101001111010001000001100100000),
            .DEVICE(DEVICE)
        )
    i_lut_590
        (
            .in_data({
                         in_data[179],
                         in_data[572],
                         in_data[553],
                         in_data[772],
                         in_data[510],
                         in_data[211]
                    }),
            .out_data(lut_590_out)
        );

reg   lut_590_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_590_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_590_ff <= lut_590_out;
    end
end

assign out_data[590] = lut_590_ff;




// LUT : 591

wire lut_591_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100000111100111111110111111110111000100100000101011110110010),
            .DEVICE(DEVICE)
        )
    i_lut_591
        (
            .in_data({
                         in_data[377],
                         in_data[196],
                         in_data[182],
                         in_data[118],
                         in_data[143],
                         in_data[420]
                    }),
            .out_data(lut_591_out)
        );

reg   lut_591_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_591_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_591_ff <= lut_591_out;
    end
end

assign out_data[591] = lut_591_ff;




// LUT : 592

wire lut_592_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110000000100000101110100011100110100000000000001101000110111),
            .DEVICE(DEVICE)
        )
    i_lut_592
        (
            .in_data({
                         in_data[695],
                         in_data[214],
                         in_data[451],
                         in_data[556],
                         in_data[586],
                         in_data[220]
                    }),
            .out_data(lut_592_out)
        );

reg   lut_592_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_592_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_592_ff <= lut_592_out;
    end
end

assign out_data[592] = lut_592_ff;




// LUT : 593

wire lut_593_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110010010101100010110010001010100000110110110100011001110000),
            .DEVICE(DEVICE)
        )
    i_lut_593
        (
            .in_data({
                         in_data[433],
                         in_data[303],
                         in_data[672],
                         in_data[629],
                         in_data[190],
                         in_data[590]
                    }),
            .out_data(lut_593_out)
        );

reg   lut_593_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_593_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_593_ff <= lut_593_out;
    end
end

assign out_data[593] = lut_593_ff;




// LUT : 594

wire lut_594_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110011011010101011101010101101101001001000001011100111110111),
            .DEVICE(DEVICE)
        )
    i_lut_594
        (
            .in_data({
                         in_data[221],
                         in_data[399],
                         in_data[782],
                         in_data[313],
                         in_data[398],
                         in_data[204]
                    }),
            .out_data(lut_594_out)
        );

reg   lut_594_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_594_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_594_ff <= lut_594_out;
    end
end

assign out_data[594] = lut_594_ff;




// LUT : 595

wire lut_595_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101001100011100010110110001110010000011000000101111111001010),
            .DEVICE(DEVICE)
        )
    i_lut_595
        (
            .in_data({
                         in_data[709],
                         in_data[348],
                         in_data[236],
                         in_data[11],
                         in_data[496],
                         in_data[294]
                    }),
            .out_data(lut_595_out)
        );

reg   lut_595_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_595_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_595_ff <= lut_595_out;
    end
end

assign out_data[595] = lut_595_ff;




// LUT : 596

wire lut_596_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010101111011100010110101011111110111100000101000110101100110),
            .DEVICE(DEVICE)
        )
    i_lut_596
        (
            .in_data({
                         in_data[32],
                         in_data[347],
                         in_data[30],
                         in_data[644],
                         in_data[517],
                         in_data[778]
                    }),
            .out_data(lut_596_out)
        );

reg   lut_596_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_596_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_596_ff <= lut_596_out;
    end
end

assign out_data[596] = lut_596_ff;




// LUT : 597

wire lut_597_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111010111001000010001000000110111010100100001101111111010100),
            .DEVICE(DEVICE)
        )
    i_lut_597
        (
            .in_data({
                         in_data[337],
                         in_data[452],
                         in_data[316],
                         in_data[387],
                         in_data[430],
                         in_data[578]
                    }),
            .out_data(lut_597_out)
        );

reg   lut_597_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_597_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_597_ff <= lut_597_out;
    end
end

assign out_data[597] = lut_597_ff;




// LUT : 598

wire lut_598_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101001010111010001010100000101010111100101011001110111100001110),
            .DEVICE(DEVICE)
        )
    i_lut_598
        (
            .in_data({
                         in_data[436],
                         in_data[36],
                         in_data[302],
                         in_data[369],
                         in_data[596],
                         in_data[127]
                    }),
            .out_data(lut_598_out)
        );

reg   lut_598_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_598_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_598_ff <= lut_598_out;
    end
end

assign out_data[598] = lut_598_ff;




// LUT : 599

wire lut_599_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110000000000101001111011000111000100001100110001111101000011),
            .DEVICE(DEVICE)
        )
    i_lut_599
        (
            .in_data({
                         in_data[150],
                         in_data[200],
                         in_data[487],
                         in_data[671],
                         in_data[187],
                         in_data[238]
                    }),
            .out_data(lut_599_out)
        );

reg   lut_599_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_599_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_599_ff <= lut_599_out;
    end
end

assign out_data[599] = lut_599_ff;




// LUT : 600

wire lut_600_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111110111000001000100010111111111001111111101110011001100),
            .DEVICE(DEVICE)
        )
    i_lut_600
        (
            .in_data({
                         in_data[343],
                         in_data[386],
                         in_data[232],
                         in_data[620],
                         in_data[354],
                         in_data[652]
                    }),
            .out_data(lut_600_out)
        );

reg   lut_600_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_600_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_600_ff <= lut_600_out;
    end
end

assign out_data[600] = lut_600_ff;




// LUT : 601

wire lut_601_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000101001001000010011000000001011100000000101111000010010101),
            .DEVICE(DEVICE)
        )
    i_lut_601
        (
            .in_data({
                         in_data[774],
                         in_data[505],
                         in_data[676],
                         in_data[781],
                         in_data[320],
                         in_data[653]
                    }),
            .out_data(lut_601_out)
        );

reg   lut_601_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_601_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_601_ff <= lut_601_out;
    end
end

assign out_data[601] = lut_601_ff;




// LUT : 602

wire lut_602_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101100111101101111001011111101100110111011011000100010101111),
            .DEVICE(DEVICE)
        )
    i_lut_602
        (
            .in_data({
                         in_data[271],
                         in_data[731],
                         in_data[222],
                         in_data[180],
                         in_data[692],
                         in_data[516]
                    }),
            .out_data(lut_602_out)
        );

reg   lut_602_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_602_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_602_ff <= lut_602_out;
    end
end

assign out_data[602] = lut_602_ff;




// LUT : 603

wire lut_603_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101110000000111010111010011001111111011111111111010100110000),
            .DEVICE(DEVICE)
        )
    i_lut_603
        (
            .in_data({
                         in_data[715],
                         in_data[603],
                         in_data[598],
                         in_data[64],
                         in_data[675],
                         in_data[237]
                    }),
            .out_data(lut_603_out)
        );

reg   lut_603_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_603_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_603_ff <= lut_603_out;
    end
end

assign out_data[603] = lut_603_ff;




// LUT : 604

wire lut_604_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101011010010110000101101000001100101010100100101111101011011),
            .DEVICE(DEVICE)
        )
    i_lut_604
        (
            .in_data({
                         in_data[685],
                         in_data[735],
                         in_data[406],
                         in_data[69],
                         in_data[270],
                         in_data[91]
                    }),
            .out_data(lut_604_out)
        );

reg   lut_604_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_604_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_604_ff <= lut_604_out;
    end
end

assign out_data[604] = lut_604_ff;




// LUT : 605

wire lut_605_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110011110000100100110010100111001010011101100000000001100110111),
            .DEVICE(DEVICE)
        )
    i_lut_605
        (
            .in_data({
                         in_data[57],
                         in_data[446],
                         in_data[693],
                         in_data[71],
                         in_data[595],
                         in_data[156]
                    }),
            .out_data(lut_605_out)
        );

reg   lut_605_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_605_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_605_ff <= lut_605_out;
    end
end

assign out_data[605] = lut_605_ff;




// LUT : 606

wire lut_606_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011011110111011011000011101101001110000101110001101001011001),
            .DEVICE(DEVICE)
        )
    i_lut_606
        (
            .in_data({
                         in_data[658],
                         in_data[284],
                         in_data[58],
                         in_data[612],
                         in_data[755],
                         in_data[459]
                    }),
            .out_data(lut_606_out)
        );

reg   lut_606_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_606_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_606_ff <= lut_606_out;
    end
end

assign out_data[606] = lut_606_ff;




// LUT : 607

wire lut_607_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010011010011111011001000100010001001100011111111101100001001),
            .DEVICE(DEVICE)
        )
    i_lut_607
        (
            .in_data({
                         in_data[634],
                         in_data[115],
                         in_data[428],
                         in_data[154],
                         in_data[260],
                         in_data[66]
                    }),
            .out_data(lut_607_out)
        );

reg   lut_607_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_607_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_607_ff <= lut_607_out;
    end
end

assign out_data[607] = lut_607_ff;




// LUT : 608

wire lut_608_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000010011100101001010110100011000011011010000001110101001001),
            .DEVICE(DEVICE)
        )
    i_lut_608
        (
            .in_data({
                         in_data[464],
                         in_data[56],
                         in_data[108],
                         in_data[231],
                         in_data[52],
                         in_data[126]
                    }),
            .out_data(lut_608_out)
        );

reg   lut_608_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_608_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_608_ff <= lut_608_out;
    end
end

assign out_data[608] = lut_608_ff;




// LUT : 609

wire lut_609_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000111000001011011110110100110110000101000001000010011000000),
            .DEVICE(DEVICE)
        )
    i_lut_609
        (
            .in_data({
                         in_data[330],
                         in_data[410],
                         in_data[257],
                         in_data[43],
                         in_data[747],
                         in_data[310]
                    }),
            .out_data(lut_609_out)
        );

reg   lut_609_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_609_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_609_ff <= lut_609_out;
    end
end

assign out_data[609] = lut_609_ff;




// LUT : 610

wire lut_610_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010010011100111110000001110110111100001111111110000101111001101),
            .DEVICE(DEVICE)
        )
    i_lut_610
        (
            .in_data({
                         in_data[152],
                         in_data[500],
                         in_data[547],
                         in_data[508],
                         in_data[605],
                         in_data[604]
                    }),
            .out_data(lut_610_out)
        );

reg   lut_610_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_610_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_610_ff <= lut_610_out;
    end
end

assign out_data[610] = lut_610_ff;




// LUT : 611

wire lut_611_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001110000111001101111001001100111011000010100101011011001101010),
            .DEVICE(DEVICE)
        )
    i_lut_611
        (
            .in_data({
                         in_data[363],
                         in_data[391],
                         in_data[323],
                         in_data[290],
                         in_data[280],
                         in_data[145]
                    }),
            .out_data(lut_611_out)
        );

reg   lut_611_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_611_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_611_ff <= lut_611_out;
    end
end

assign out_data[611] = lut_611_ff;




// LUT : 612

wire lut_612_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101111001001011100110011111110111100011100000111000001110000),
            .DEVICE(DEVICE)
        )
    i_lut_612
        (
            .in_data({
                         in_data[48],
                         in_data[581],
                         in_data[184],
                         in_data[131],
                         in_data[140],
                         in_data[512]
                    }),
            .out_data(lut_612_out)
        );

reg   lut_612_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_612_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_612_ff <= lut_612_out;
    end
end

assign out_data[612] = lut_612_ff;




// LUT : 613

wire lut_613_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110110010101100101000000111100001010110100101101011000100001100),
            .DEVICE(DEVICE)
        )
    i_lut_613
        (
            .in_data({
                         in_data[424],
                         in_data[219],
                         in_data[607],
                         in_data[616],
                         in_data[750],
                         in_data[515]
                    }),
            .out_data(lut_613_out)
        );

reg   lut_613_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_613_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_613_ff <= lut_613_out;
    end
end

assign out_data[613] = lut_613_ff;




// LUT : 614

wire lut_614_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000000111000101001110101110100000110011011101110101100010000),
            .DEVICE(DEVICE)
        )
    i_lut_614
        (
            .in_data({
                         in_data[248],
                         in_data[783],
                         in_data[307],
                         in_data[627],
                         in_data[25],
                         in_data[382]
                    }),
            .out_data(lut_614_out)
        );

reg   lut_614_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_614_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_614_ff <= lut_614_out;
    end
end

assign out_data[614] = lut_614_ff;




// LUT : 615

wire lut_615_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110101011110000010010001110000101110111110101100100010001001111),
            .DEVICE(DEVICE)
        )
    i_lut_615
        (
            .in_data({
                         in_data[403],
                         in_data[765],
                         in_data[522],
                         in_data[375],
                         in_data[312],
                         in_data[82]
                    }),
            .out_data(lut_615_out)
        );

reg   lut_615_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_615_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_615_ff <= lut_615_out;
    end
end

assign out_data[615] = lut_615_ff;




// LUT : 616

wire lut_616_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100000010011110000000001010110001000000100100010111010101001),
            .DEVICE(DEVICE)
        )
    i_lut_616
        (
            .in_data({
                         in_data[437],
                         in_data[288],
                         in_data[163],
                         in_data[341],
                         in_data[758],
                         in_data[727]
                    }),
            .out_data(lut_616_out)
        );

reg   lut_616_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_616_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_616_ff <= lut_616_out;
    end
end

assign out_data[616] = lut_616_ff;




// LUT : 617

wire lut_617_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001110000101001110010110011100011100111110001110000111101110000),
            .DEVICE(DEVICE)
        )
    i_lut_617
        (
            .in_data({
                         in_data[471],
                         in_data[34],
                         in_data[159],
                         in_data[0],
                         in_data[647],
                         in_data[746]
                    }),
            .out_data(lut_617_out)
        );

reg   lut_617_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_617_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_617_ff <= lut_617_out;
    end
end

assign out_data[617] = lut_617_ff;




// LUT : 618

wire lut_618_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101001110111011000001100011100011110110100110100000011001111),
            .DEVICE(DEVICE)
        )
    i_lut_618
        (
            .in_data({
                         in_data[599],
                         in_data[335],
                         in_data[16],
                         in_data[175],
                         in_data[134],
                         in_data[304]
                    }),
            .out_data(lut_618_out)
        );

reg   lut_618_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_618_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_618_ff <= lut_618_out;
    end
end

assign out_data[618] = lut_618_ff;




// LUT : 619

wire lut_619_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010110110100001111010011101011010001100000110100101000001011),
            .DEVICE(DEVICE)
        )
    i_lut_619
        (
            .in_data({
                         in_data[26],
                         in_data[149],
                         in_data[421],
                         in_data[315],
                         in_data[681],
                         in_data[732]
                    }),
            .out_data(lut_619_out)
        );

reg   lut_619_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_619_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_619_ff <= lut_619_out;
    end
end

assign out_data[619] = lut_619_ff;




// LUT : 620

wire lut_620_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001011010100100000110001010000111010010110111100011100000001101),
            .DEVICE(DEVICE)
        )
    i_lut_620
        (
            .in_data({
                         in_data[98],
                         in_data[144],
                         in_data[762],
                         in_data[78],
                         in_data[356],
                         in_data[716]
                    }),
            .out_data(lut_620_out)
        );

reg   lut_620_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_620_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_620_ff <= lut_620_out;
    end
end

assign out_data[620] = lut_620_ff;




// LUT : 621

wire lut_621_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100111101010001101110111011111001011011100001011101111011101),
            .DEVICE(DEVICE)
        )
    i_lut_621
        (
            .in_data({
                         in_data[367],
                         in_data[361],
                         in_data[394],
                         in_data[463],
                         in_data[192],
                         in_data[245]
                    }),
            .out_data(lut_621_out)
        );

reg   lut_621_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_621_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_621_ff <= lut_621_out;
    end
end

assign out_data[621] = lut_621_ff;




// LUT : 622

wire lut_622_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000111011001101010011001000001111000111001011100010001000101),
            .DEVICE(DEVICE)
        )
    i_lut_622
        (
            .in_data({
                         in_data[106],
                         in_data[654],
                         in_data[185],
                         in_data[223],
                         in_data[254],
                         in_data[568]
                    }),
            .out_data(lut_622_out)
        );

reg   lut_622_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_622_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_622_ff <= lut_622_out;
    end
end

assign out_data[622] = lut_622_ff;




// LUT : 623

wire lut_623_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000100000101001001000011100000010001100010000010001000101100111),
            .DEVICE(DEVICE)
        )
    i_lut_623
        (
            .in_data({
                         in_data[47],
                         in_data[178],
                         in_data[389],
                         in_data[626],
                         in_data[6],
                         in_data[472]
                    }),
            .out_data(lut_623_out)
        );

reg   lut_623_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_623_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_623_ff <= lut_623_out;
    end
end

assign out_data[623] = lut_623_ff;




// LUT : 624

wire lut_624_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101000110001101110100111100101000100001111110100111001111110),
            .DEVICE(DEVICE)
        )
    i_lut_624
        (
            .in_data({
                         in_data[28],
                         in_data[743],
                         in_data[587],
                         in_data[560],
                         in_data[283],
                         in_data[287]
                    }),
            .out_data(lut_624_out)
        );

reg   lut_624_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_624_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_624_ff <= lut_624_out;
    end
end

assign out_data[624] = lut_624_ff;




// LUT : 625

wire lut_625_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101111101011101111101101001100110111010101101000110011001010),
            .DEVICE(DEVICE)
        )
    i_lut_625
        (
            .in_data({
                         in_data[86],
                         in_data[588],
                         in_data[773],
                         in_data[691],
                         in_data[210],
                         in_data[539]
                    }),
            .out_data(lut_625_out)
        );

reg   lut_625_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_625_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_625_ff <= lut_625_out;
    end
end

assign out_data[625] = lut_625_ff;




// LUT : 626

wire lut_626_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100011001110111000001011001011111011110110111000010001000000000),
            .DEVICE(DEVICE)
        )
    i_lut_626
        (
            .in_data({
                         in_data[42],
                         in_data[366],
                         in_data[325],
                         in_data[585],
                         in_data[666],
                         in_data[650]
                    }),
            .out_data(lut_626_out)
        );

reg   lut_626_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_626_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_626_ff <= lut_626_out;
    end
end

assign out_data[626] = lut_626_ff;




// LUT : 627

wire lut_627_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001111111000011001001111100111101101001000110011010011100100010),
            .DEVICE(DEVICE)
        )
    i_lut_627
        (
            .in_data({
                         in_data[105],
                         in_data[170],
                         in_data[174],
                         in_data[645],
                         in_data[729],
                         in_data[648]
                    }),
            .out_data(lut_627_out)
        );

reg   lut_627_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_627_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_627_ff <= lut_627_out;
    end
end

assign out_data[627] = lut_627_ff;




// LUT : 628

wire lut_628_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000011110010011100011001101110001100111000111111110110111011100),
            .DEVICE(DEVICE)
        )
    i_lut_628
        (
            .in_data({
                         in_data[216],
                         in_data[75],
                         in_data[442],
                         in_data[611],
                         in_data[90],
                         in_data[258]
                    }),
            .out_data(lut_628_out)
        );

reg   lut_628_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_628_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_628_ff <= lut_628_out;
    end
end

assign out_data[628] = lut_628_ff;




// LUT : 629

wire lut_629_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100001001100100100101001010001110000101011101111000011100001),
            .DEVICE(DEVICE)
        )
    i_lut_629
        (
            .in_data({
                         in_data[478],
                         in_data[365],
                         in_data[132],
                         in_data[89],
                         in_data[413],
                         in_data[523]
                    }),
            .out_data(lut_629_out)
        );

reg   lut_629_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_629_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_629_ff <= lut_629_out;
    end
end

assign out_data[629] = lut_629_ff;




// LUT : 630

wire lut_630_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111111111111111000111111111101001100011011001111011111001100),
            .DEVICE(DEVICE)
        )
    i_lut_630
        (
            .in_data({
                         in_data[195],
                         in_data[193],
                         in_data[116],
                         in_data[267],
                         in_data[171],
                         in_data[520]
                    }),
            .out_data(lut_630_out)
        );

reg   lut_630_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_630_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_630_ff <= lut_630_out;
    end
end

assign out_data[630] = lut_630_ff;




// LUT : 631

wire lut_631_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111101110101111111111011111101010011111111010111011110111111),
            .DEVICE(DEVICE)
        )
    i_lut_631
        (
            .in_data({
                         in_data[234],
                         in_data[637],
                         in_data[651],
                         in_data[226],
                         in_data[481],
                         in_data[631]
                    }),
            .out_data(lut_631_out)
        );

reg   lut_631_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_631_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_631_ff <= lut_631_out;
    end
end

assign out_data[631] = lut_631_ff;




// LUT : 632

wire lut_632_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010100010010011001011101000100010010010001100000110001100110),
            .DEVICE(DEVICE)
        )
    i_lut_632
        (
            .in_data({
                         in_data[748],
                         in_data[609],
                         in_data[411],
                         in_data[711],
                         in_data[706],
                         in_data[137]
                    }),
            .out_data(lut_632_out)
        );

reg   lut_632_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_632_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_632_ff <= lut_632_out;
    end
end

assign out_data[632] = lut_632_ff;




// LUT : 633

wire lut_633_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001000100011111111111011001000110010100101011111111100001100),
            .DEVICE(DEVICE)
        )
    i_lut_633
        (
            .in_data({
                         in_data[77],
                         in_data[33],
                         in_data[484],
                         in_data[649],
                         in_data[613],
                         in_data[129]
                    }),
            .out_data(lut_633_out)
        );

reg   lut_633_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_633_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_633_ff <= lut_633_out;
    end
end

assign out_data[633] = lut_633_ff;




// LUT : 634

wire lut_634_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100000110000110001010000010000101011010101011010000111111001),
            .DEVICE(DEVICE)
        )
    i_lut_634
        (
            .in_data({
                         in_data[164],
                         in_data[660],
                         in_data[432],
                         in_data[201],
                         in_data[111],
                         in_data[526]
                    }),
            .out_data(lut_634_out)
        );

reg   lut_634_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_634_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_634_ff <= lut_634_out;
    end
end

assign out_data[634] = lut_634_ff;




// LUT : 635

wire lut_635_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111100111111001100101110101000011011000111110011101010101010),
            .DEVICE(DEVICE)
        )
    i_lut_635
        (
            .in_data({
                         in_data[665],
                         in_data[266],
                         in_data[165],
                         in_data[191],
                         in_data[117],
                         in_data[125]
                    }),
            .out_data(lut_635_out)
        );

reg   lut_635_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_635_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_635_ff <= lut_635_out;
    end
end

assign out_data[635] = lut_635_ff;




// LUT : 636

wire lut_636_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010100101110010001010001011010000011001000010110000001000000),
            .DEVICE(DEVICE)
        )
    i_lut_636
        (
            .in_data({
                         in_data[35],
                         in_data[276],
                         in_data[677],
                         in_data[564],
                         in_data[737],
                         in_data[1]
                    }),
            .out_data(lut_636_out)
        );

reg   lut_636_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_636_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_636_ff <= lut_636_out;
    end
end

assign out_data[636] = lut_636_ff;




// LUT : 637

wire lut_637_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001100101010101011100011011010101111101100110001011110110110010),
            .DEVICE(DEVICE)
        )
    i_lut_637
        (
            .in_data({
                         in_data[110],
                         in_data[456],
                         in_data[624],
                         in_data[239],
                         in_data[10],
                         in_data[469]
                    }),
            .out_data(lut_637_out)
        );

reg   lut_637_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_637_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_637_ff <= lut_637_out;
    end
end

assign out_data[637] = lut_637_ff;




// LUT : 638

wire lut_638_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110010011010110111100111111011101000111000111010111110000000),
            .DEVICE(DEVICE)
        )
    i_lut_638
        (
            .in_data({
                         in_data[431],
                         in_data[87],
                         in_data[202],
                         in_data[717],
                         in_data[409],
                         in_data[72]
                    }),
            .out_data(lut_638_out)
        );

reg   lut_638_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_638_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_638_ff <= lut_638_out;
    end
end

assign out_data[638] = lut_638_ff;




// LUT : 639

wire lut_639_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001011001100111010000000000011010100000000000001011100000011),
            .DEVICE(DEVICE)
        )
    i_lut_639
        (
            .in_data({
                         in_data[779],
                         in_data[721],
                         in_data[8],
                         in_data[427],
                         in_data[282],
                         in_data[256]
                    }),
            .out_data(lut_639_out)
        );

reg   lut_639_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_639_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_639_ff <= lut_639_out;
    end
end

assign out_data[639] = lut_639_ff;




// LUT : 640

wire lut_640_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001001011011111011011111000000100111111110101000010100000010),
            .DEVICE(DEVICE)
        )
    i_lut_640
        (
            .in_data({
                         in_data[720],
                         in_data[618],
                         in_data[61],
                         in_data[103],
                         in_data[352],
                         in_data[251]
                    }),
            .out_data(lut_640_out)
        );

reg   lut_640_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_640_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_640_ff <= lut_640_out;
    end
end

assign out_data[640] = lut_640_ff;




// LUT : 641

wire lut_641_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101001110011010000010001100111111111111111111111111011101010),
            .DEVICE(DEVICE)
        )
    i_lut_641
        (
            .in_data({
                         in_data[726],
                         in_data[93],
                         in_data[511],
                         in_data[554],
                         in_data[181],
                         in_data[158]
                    }),
            .out_data(lut_641_out)
        );

reg   lut_641_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_641_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_641_ff <= lut_641_out;
    end
end

assign out_data[641] = lut_641_ff;




// LUT : 642

wire lut_642_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000010100101000000000000010000110011000000110100011100000111),
            .DEVICE(DEVICE)
        )
    i_lut_642
        (
            .in_data({
                         in_data[659],
                         in_data[480],
                         in_data[486],
                         in_data[576],
                         in_data[630],
                         in_data[319]
                    }),
            .out_data(lut_642_out)
        );

reg   lut_642_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_642_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_642_ff <= lut_642_out;
    end
end

assign out_data[642] = lut_642_ff;




// LUT : 643

wire lut_643_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010010011010011000001010101111001111011011110011000111001111110),
            .DEVICE(DEVICE)
        )
    i_lut_643
        (
            .in_data({
                         in_data[507],
                         in_data[532],
                         in_data[228],
                         in_data[55],
                         in_data[124],
                         in_data[655]
                    }),
            .out_data(lut_643_out)
        );

reg   lut_643_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_643_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_643_ff <= lut_643_out;
    end
end

assign out_data[643] = lut_643_ff;




// LUT : 644

wire lut_644_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000100010011110110010011111100011101110111111010000011001100),
            .DEVICE(DEVICE)
        )
    i_lut_644
        (
            .in_data({
                         in_data[619],
                         in_data[104],
                         in_data[759],
                         in_data[328],
                         in_data[74],
                         in_data[289]
                    }),
            .out_data(lut_644_out)
        );

reg   lut_644_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_644_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_644_ff <= lut_644_out;
    end
end

assign out_data[644] = lut_644_ff;




// LUT : 645

wire lut_645_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010001101100000001000100010010000000001111110000101000000000),
            .DEVICE(DEVICE)
        )
    i_lut_645
        (
            .in_data({
                         in_data[97],
                         in_data[274],
                         in_data[535],
                         in_data[602],
                         in_data[80],
                         in_data[208]
                    }),
            .out_data(lut_645_out)
        );

reg   lut_645_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_645_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_645_ff <= lut_645_out;
    end
end

assign out_data[645] = lut_645_ff;




// LUT : 646

wire lut_646_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000010011010000011001010100010000111100000100101110111101111),
            .DEVICE(DEVICE)
        )
    i_lut_646
        (
            .in_data({
                         in_data[83],
                         in_data[518],
                         in_data[503],
                         in_data[344],
                         in_data[101],
                         in_data[24]
                    }),
            .out_data(lut_646_out)
        );

reg   lut_646_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_646_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_646_ff <= lut_646_out;
    end
end

assign out_data[646] = lut_646_ff;




// LUT : 647

wire lut_647_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111011110110110001111000101000001100111100001111110010011100),
            .DEVICE(DEVICE)
        )
    i_lut_647
        (
            .in_data({
                         in_data[763],
                         in_data[416],
                         in_data[661],
                         in_data[139],
                         in_data[141],
                         in_data[610]
                    }),
            .out_data(lut_647_out)
        );

reg   lut_647_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_647_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_647_ff <= lut_647_out;
    end
end

assign out_data[647] = lut_647_ff;




// LUT : 648

wire lut_648_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100101010001010000010010000000110001010110010010100100100000),
            .DEVICE(DEVICE)
        )
    i_lut_648
        (
            .in_data({
                         in_data[570],
                         in_data[286],
                         in_data[571],
                         in_data[447],
                         in_data[592],
                         in_data[668]
                    }),
            .out_data(lut_648_out)
        );

reg   lut_648_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_648_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_648_ff <= lut_648_out;
    end
end

assign out_data[648] = lut_648_ff;




// LUT : 649

wire lut_649_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000011001011111100000100001100011110110011111011111101000011),
            .DEVICE(DEVICE)
        )
    i_lut_649
        (
            .in_data({
                         in_data[233],
                         in_data[355],
                         in_data[29],
                         in_data[577],
                         in_data[769],
                         in_data[397]
                    }),
            .out_data(lut_649_out)
        );

reg   lut_649_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_649_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_649_ff <= lut_649_out;
    end
end

assign out_data[649] = lut_649_ff;




// LUT : 650

wire lut_650_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100001110100010010010011010000001111111011110000101100111001000),
            .DEVICE(DEVICE)
        )
    i_lut_650
        (
            .in_data({
                         in_data[232],
                         in_data[518],
                         in_data[20],
                         in_data[670],
                         in_data[265],
                         in_data[19]
                    }),
            .out_data(lut_650_out)
        );

reg   lut_650_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_650_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_650_ff <= lut_650_out;
    end
end

assign out_data[650] = lut_650_ff;




// LUT : 651

wire lut_651_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001011100100000001101000000000000111110000000000011110100),
            .DEVICE(DEVICE)
        )
    i_lut_651
        (
            .in_data({
                         in_data[695],
                         in_data[625],
                         in_data[634],
                         in_data[709],
                         in_data[267],
                         in_data[597]
                    }),
            .out_data(lut_651_out)
        );

reg   lut_651_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_651_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_651_ff <= lut_651_out;
    end
end

assign out_data[651] = lut_651_ff;




// LUT : 652

wire lut_652_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010000101111111111111111111100101010111001001110111011110100),
            .DEVICE(DEVICE)
        )
    i_lut_652
        (
            .in_data({
                         in_data[495],
                         in_data[641],
                         in_data[575],
                         in_data[456],
                         in_data[494],
                         in_data[42]
                    }),
            .out_data(lut_652_out)
        );

reg   lut_652_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_652_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_652_ff <= lut_652_out;
    end
end

assign out_data[652] = lut_652_ff;




// LUT : 653

wire lut_653_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001011100011101111000001110010110111111011110110011101101101011),
            .DEVICE(DEVICE)
        )
    i_lut_653
        (
            .in_data({
                         in_data[770],
                         in_data[154],
                         in_data[524],
                         in_data[4],
                         in_data[437],
                         in_data[256]
                    }),
            .out_data(lut_653_out)
        );

reg   lut_653_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_653_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_653_ff <= lut_653_out;
    end
end

assign out_data[653] = lut_653_ff;




// LUT : 654

wire lut_654_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000001100000010100001111010010110101011111110001000000101111),
            .DEVICE(DEVICE)
        )
    i_lut_654
        (
            .in_data({
                         in_data[512],
                         in_data[647],
                         in_data[301],
                         in_data[731],
                         in_data[204],
                         in_data[608]
                    }),
            .out_data(lut_654_out)
        );

reg   lut_654_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_654_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_654_ff <= lut_654_out;
    end
end

assign out_data[654] = lut_654_ff;




// LUT : 655

wire lut_655_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000011000100100110010010001100100010101011100010000110000010101),
            .DEVICE(DEVICE)
        )
    i_lut_655
        (
            .in_data({
                         in_data[773],
                         in_data[728],
                         in_data[213],
                         in_data[183],
                         in_data[149],
                         in_data[122]
                    }),
            .out_data(lut_655_out)
        );

reg   lut_655_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_655_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_655_ff <= lut_655_out;
    end
end

assign out_data[655] = lut_655_ff;




// LUT : 656

wire lut_656_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111101111101101101111011110100111101011111010101100110111100),
            .DEVICE(DEVICE)
        )
    i_lut_656
        (
            .in_data({
                         in_data[384],
                         in_data[548],
                         in_data[352],
                         in_data[94],
                         in_data[422],
                         in_data[545]
                    }),
            .out_data(lut_656_out)
        );

reg   lut_656_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_656_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_656_ff <= lut_656_out;
    end
end

assign out_data[656] = lut_656_ff;




// LUT : 657

wire lut_657_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001100000010011011100011111111100000100000001100010001100100111),
            .DEVICE(DEVICE)
        )
    i_lut_657
        (
            .in_data({
                         in_data[145],
                         in_data[473],
                         in_data[315],
                         in_data[292],
                         in_data[656],
                         in_data[637]
                    }),
            .out_data(lut_657_out)
        );

reg   lut_657_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_657_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_657_ff <= lut_657_out;
    end
end

assign out_data[657] = lut_657_ff;




// LUT : 658

wire lut_658_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001000000100011110100101100110011000001011101101110010000101),
            .DEVICE(DEVICE)
        )
    i_lut_658
        (
            .in_data({
                         in_data[513],
                         in_data[452],
                         in_data[326],
                         in_data[50],
                         in_data[110],
                         in_data[13]
                    }),
            .out_data(lut_658_out)
        );

reg   lut_658_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_658_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_658_ff <= lut_658_out;
    end
end

assign out_data[658] = lut_658_ff;




// LUT : 659

wire lut_659_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110110110000000010100100000111101110111010101010000100011000101),
            .DEVICE(DEVICE)
        )
    i_lut_659
        (
            .in_data({
                         in_data[203],
                         in_data[115],
                         in_data[138],
                         in_data[603],
                         in_data[133],
                         in_data[393]
                    }),
            .out_data(lut_659_out)
        );

reg   lut_659_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_659_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_659_ff <= lut_659_out;
    end
end

assign out_data[659] = lut_659_ff;




// LUT : 660

wire lut_660_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100011011110111010011011111111111100001101110000111001010111010),
            .DEVICE(DEVICE)
        )
    i_lut_660
        (
            .in_data({
                         in_data[611],
                         in_data[275],
                         in_data[17],
                         in_data[537],
                         in_data[485],
                         in_data[638]
                    }),
            .out_data(lut_660_out)
        );

reg   lut_660_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_660_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_660_ff <= lut_660_out;
    end
end

assign out_data[660] = lut_660_ff;




// LUT : 661

wire lut_661_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000011110011000011011001011101100110110001000000010000000001111),
            .DEVICE(DEVICE)
        )
    i_lut_661
        (
            .in_data({
                         in_data[8],
                         in_data[226],
                         in_data[617],
                         in_data[642],
                         in_data[233],
                         in_data[380]
                    }),
            .out_data(lut_661_out)
        );

reg   lut_661_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_661_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_661_ff <= lut_661_out;
    end
end

assign out_data[661] = lut_661_ff;




// LUT : 662

wire lut_662_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000100110100000000111010001100011101100100001010000000000111100),
            .DEVICE(DEVICE)
        )
    i_lut_662
        (
            .in_data({
                         in_data[58],
                         in_data[211],
                         in_data[108],
                         in_data[766],
                         in_data[706],
                         in_data[102]
                    }),
            .out_data(lut_662_out)
        );

reg   lut_662_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_662_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_662_ff <= lut_662_out;
    end
end

assign out_data[662] = lut_662_ff;




// LUT : 663

wire lut_663_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101000101010100111110001100100001000011001010011100100010001),
            .DEVICE(DEVICE)
        )
    i_lut_663
        (
            .in_data({
                         in_data[397],
                         in_data[509],
                         in_data[755],
                         in_data[97],
                         in_data[475],
                         in_data[46]
                    }),
            .out_data(lut_663_out)
        );

reg   lut_663_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_663_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_663_ff <= lut_663_out;
    end
end

assign out_data[663] = lut_663_ff;




// LUT : 664

wire lut_664_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111001010000100011000100010010000110110101001010100101010000100),
            .DEVICE(DEVICE)
        )
    i_lut_664
        (
            .in_data({
                         in_data[543],
                         in_data[493],
                         in_data[26],
                         in_data[36],
                         in_data[436],
                         in_data[746]
                    }),
            .out_data(lut_664_out)
        );

reg   lut_664_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_664_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_664_ff <= lut_664_out;
    end
end

assign out_data[664] = lut_664_ff;




// LUT : 665

wire lut_665_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100110100111101000001110101011111110000000011011000111000100),
            .DEVICE(DEVICE)
        )
    i_lut_665
        (
            .in_data({
                         in_data[663],
                         in_data[182],
                         in_data[27],
                         in_data[168],
                         in_data[399],
                         in_data[31]
                    }),
            .out_data(lut_665_out)
        );

reg   lut_665_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_665_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_665_ff <= lut_665_out;
    end
end

assign out_data[665] = lut_665_ff;




// LUT : 666

wire lut_666_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000010010101000110101110010100100101001001000111111101110000),
            .DEVICE(DEVICE)
        )
    i_lut_666
        (
            .in_data({
                         in_data[314],
                         in_data[579],
                         in_data[254],
                         in_data[503],
                         in_data[287],
                         in_data[407]
                    }),
            .out_data(lut_666_out)
        );

reg   lut_666_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_666_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_666_ff <= lut_666_out;
    end
end

assign out_data[666] = lut_666_ff;




// LUT : 667

wire lut_667_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010010101000010110100010100011010000000010001111000011100000),
            .DEVICE(DEVICE)
        )
    i_lut_667
        (
            .in_data({
                         in_data[239],
                         in_data[426],
                         in_data[609],
                         in_data[570],
                         in_data[351],
                         in_data[588]
                    }),
            .out_data(lut_667_out)
        );

reg   lut_667_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_667_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_667_ff <= lut_667_out;
    end
end

assign out_data[667] = lut_667_ff;




// LUT : 668

wire lut_668_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101001110000000001000000110011100111101010010011111011100001010),
            .DEVICE(DEVICE)
        )
    i_lut_668
        (
            .in_data({
                         in_data[289],
                         in_data[139],
                         in_data[771],
                         in_data[0],
                         in_data[685],
                         in_data[750]
                    }),
            .out_data(lut_668_out)
        );

reg   lut_668_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_668_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_668_ff <= lut_668_out;
    end
end

assign out_data[668] = lut_668_ff;




// LUT : 669

wire lut_669_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000001110000000111001110110101010110111111110111110010111111),
            .DEVICE(DEVICE)
        )
    i_lut_669
        (
            .in_data({
                         in_data[521],
                         in_data[623],
                         in_data[159],
                         in_data[740],
                         in_data[76],
                         in_data[405]
                    }),
            .out_data(lut_669_out)
        );

reg   lut_669_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_669_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_669_ff <= lut_669_out;
    end
end

assign out_data[669] = lut_669_ff;




// LUT : 670

wire lut_670_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000101100111000000110101101001101010100001111101010111011100),
            .DEVICE(DEVICE)
        )
    i_lut_670
        (
            .in_data({
                         in_data[774],
                         in_data[699],
                         in_data[569],
                         in_data[334],
                         in_data[360],
                         in_data[74]
                    }),
            .out_data(lut_670_out)
        );

reg   lut_670_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_670_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_670_ff <= lut_670_out;
    end
end

assign out_data[670] = lut_670_ff;




// LUT : 671

wire lut_671_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101001001111011000101110011101101111001001100111110110110001000),
            .DEVICE(DEVICE)
        )
    i_lut_671
        (
            .in_data({
                         in_data[250],
                         in_data[359],
                         in_data[80],
                         in_data[630],
                         in_data[170],
                         in_data[259]
                    }),
            .out_data(lut_671_out)
        );

reg   lut_671_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_671_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_671_ff <= lut_671_out;
    end
end

assign out_data[671] = lut_671_ff;




// LUT : 672

wire lut_672_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111010011101000110001101110111111010101011100101101111011100),
            .DEVICE(DEVICE)
        )
    i_lut_672
        (
            .in_data({
                         in_data[269],
                         in_data[82],
                         in_data[756],
                         in_data[566],
                         in_data[332],
                         in_data[161]
                    }),
            .out_data(lut_672_out)
        );

reg   lut_672_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_672_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_672_ff <= lut_672_out;
    end
end

assign out_data[672] = lut_672_ff;




// LUT : 673

wire lut_673_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111001000011011010001010110100010010111000100011000011010111100),
            .DEVICE(DEVICE)
        )
    i_lut_673
        (
            .in_data({
                         in_data[615],
                         in_data[209],
                         in_data[451],
                         in_data[747],
                         in_data[729],
                         in_data[419]
                    }),
            .out_data(lut_673_out)
        );

reg   lut_673_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_673_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_673_ff <= lut_673_out;
    end
end

assign out_data[673] = lut_673_ff;




// LUT : 674

wire lut_674_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111000100011000011111111111010111001101100111010111011111010),
            .DEVICE(DEVICE)
        )
    i_lut_674
        (
            .in_data({
                         in_data[539],
                         in_data[767],
                         in_data[660],
                         in_data[574],
                         in_data[175],
                         in_data[236]
                    }),
            .out_data(lut_674_out)
        );

reg   lut_674_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_674_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_674_ff <= lut_674_out;
    end
end

assign out_data[674] = lut_674_ff;




// LUT : 675

wire lut_675_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011110110010100000001011100100100110011010000000010000000000),
            .DEVICE(DEVICE)
        )
    i_lut_675
        (
            .in_data({
                         in_data[458],
                         in_data[689],
                         in_data[64],
                         in_data[434],
                         in_data[646],
                         in_data[578]
                    }),
            .out_data(lut_675_out)
        );

reg   lut_675_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_675_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_675_ff <= lut_675_out;
    end
end

assign out_data[675] = lut_675_ff;




// LUT : 676

wire lut_676_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110110001101011010101000001000010110011100011111011010010100110),
            .DEVICE(DEVICE)
        )
    i_lut_676
        (
            .in_data({
                         in_data[704],
                         in_data[697],
                         in_data[542],
                         in_data[590],
                         in_data[123],
                         in_data[375]
                    }),
            .out_data(lut_676_out)
        );

reg   lut_676_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_676_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_676_ff <= lut_676_out;
    end
end

assign out_data[676] = lut_676_ff;




// LUT : 677

wire lut_677_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100110000000001100001011100001011001111111001010000001000001),
            .DEVICE(DEVICE)
        )
    i_lut_677
        (
            .in_data({
                         in_data[44],
                         in_data[144],
                         in_data[156],
                         in_data[640],
                         in_data[438],
                         in_data[716]
                    }),
            .out_data(lut_677_out)
        );

reg   lut_677_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_677_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_677_ff <= lut_677_out;
    end
end

assign out_data[677] = lut_677_ff;




// LUT : 678

wire lut_678_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110101101001111011000010110001101100111010000010011000110011),
            .DEVICE(DEVICE)
        )
    i_lut_678
        (
            .in_data({
                         in_data[772],
                         in_data[51],
                         in_data[143],
                         in_data[317],
                         in_data[506],
                         in_data[340]
                    }),
            .out_data(lut_678_out)
        );

reg   lut_678_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_678_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_678_ff <= lut_678_out;
    end
end

assign out_data[678] = lut_678_ff;




// LUT : 679

wire lut_679_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110101000101100000101010000110110111101111110001011101000010010),
            .DEVICE(DEVICE)
        )
    i_lut_679
        (
            .in_data({
                         in_data[169],
                         in_data[576],
                         in_data[52],
                         in_data[477],
                         in_data[33],
                         in_data[761]
                    }),
            .out_data(lut_679_out)
        );

reg   lut_679_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_679_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_679_ff <= lut_679_out;
    end
end

assign out_data[679] = lut_679_ff;




// LUT : 680

wire lut_680_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001001111111101011111111010000010001010000010001010111000001),
            .DEVICE(DEVICE)
        )
    i_lut_680
        (
            .in_data({
                         in_data[418],
                         in_data[550],
                         in_data[202],
                         in_data[564],
                         in_data[769],
                         in_data[207]
                    }),
            .out_data(lut_680_out)
        );

reg   lut_680_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_680_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_680_ff <= lut_680_out;
    end
end

assign out_data[680] = lut_680_ff;




// LUT : 681

wire lut_681_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000100010111011110111001011101001101100010111010011110010),
            .DEVICE(DEVICE)
        )
    i_lut_681
        (
            .in_data({
                         in_data[627],
                         in_data[273],
                         in_data[147],
                         in_data[179],
                         in_data[111],
                         in_data[691]
                    }),
            .out_data(lut_681_out)
        );

reg   lut_681_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_681_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_681_ff <= lut_681_out;
    end
end

assign out_data[681] = lut_681_ff;




// LUT : 682

wire lut_682_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010110100101010000100011111111100011101111110000101011110011),
            .DEVICE(DEVICE)
        )
    i_lut_682
        (
            .in_data({
                         in_data[748],
                         in_data[727],
                         in_data[469],
                         in_data[215],
                         in_data[343],
                         in_data[324]
                    }),
            .out_data(lut_682_out)
        );

reg   lut_682_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_682_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_682_ff <= lut_682_out;
    end
end

assign out_data[682] = lut_682_ff;




// LUT : 683

wire lut_683_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010001001000100100111010100101011110000010100010010100010001),
            .DEVICE(DEVICE)
        )
    i_lut_683
        (
            .in_data({
                         in_data[37],
                         in_data[53],
                         in_data[246],
                         in_data[768],
                         in_data[140],
                         in_data[679]
                    }),
            .out_data(lut_683_out)
        );

reg   lut_683_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_683_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_683_ff <= lut_683_out;
    end
end

assign out_data[683] = lut_683_ff;




// LUT : 684

wire lut_684_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111111001010111000110110101111100100111101111100110111001101),
            .DEVICE(DEVICE)
        )
    i_lut_684
        (
            .in_data({
                         in_data[196],
                         in_data[459],
                         in_data[629],
                         in_data[303],
                         in_data[228],
                         in_data[356]
                    }),
            .out_data(lut_684_out)
        );

reg   lut_684_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_684_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_684_ff <= lut_684_out;
    end
end

assign out_data[684] = lut_684_ff;




// LUT : 685

wire lut_685_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001011100010000000010011001100000001110001000010011100100011),
            .DEVICE(DEVICE)
        )
    i_lut_685
        (
            .in_data({
                         in_data[187],
                         in_data[555],
                         in_data[462],
                         in_data[567],
                         in_data[105],
                         in_data[398]
                    }),
            .out_data(lut_685_out)
        );

reg   lut_685_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_685_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_685_ff <= lut_685_out;
    end
end

assign out_data[685] = lut_685_ff;




// LUT : 686

wire lut_686_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110001001000100010000110100111111000001010000111011011101001),
            .DEVICE(DEVICE)
        )
    i_lut_686
        (
            .in_data({
                         in_data[491],
                         in_data[723],
                         in_data[502],
                         in_data[667],
                         in_data[79],
                         in_data[676]
                    }),
            .out_data(lut_686_out)
        );

reg   lut_686_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_686_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_686_ff <= lut_686_out;
    end
end

assign out_data[686] = lut_686_ff;




// LUT : 687

wire lut_687_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001010001000101110111110001101101110110001111111010001111111),
            .DEVICE(DEVICE)
        )
    i_lut_687
        (
            .in_data({
                         in_data[732],
                         in_data[21],
                         in_data[406],
                         in_data[253],
                         in_data[738],
                         in_data[258]
                    }),
            .out_data(lut_687_out)
        );

reg   lut_687_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_687_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_687_ff <= lut_687_out;
    end
end

assign out_data[687] = lut_687_ff;




// LUT : 688

wire lut_688_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101110011100011001111101100001110110000000011010011110110011),
            .DEVICE(DEVICE)
        )
    i_lut_688
        (
            .in_data({
                         in_data[9],
                         in_data[528],
                         in_data[562],
                         in_data[220],
                         in_data[572],
                         in_data[514]
                    }),
            .out_data(lut_688_out)
        );

reg   lut_688_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_688_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_688_ff <= lut_688_out;
    end
end

assign out_data[688] = lut_688_ff;




// LUT : 689

wire lut_689_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001100111001101001111001000000110100010000110110000111001000111),
            .DEVICE(DEVICE)
        )
    i_lut_689
        (
            .in_data({
                         in_data[632],
                         in_data[77],
                         in_data[613],
                         in_data[450],
                         in_data[70],
                         in_data[229]
                    }),
            .out_data(lut_689_out)
        );

reg   lut_689_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_689_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_689_ff <= lut_689_out;
    end
end

assign out_data[689] = lut_689_ff;




// LUT : 690

wire lut_690_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101010011010011111011011001001110011010110100111111110011010),
            .DEVICE(DEVICE)
        )
    i_lut_690
        (
            .in_data({
                         in_data[775],
                         in_data[271],
                         in_data[176],
                         in_data[63],
                         in_data[776],
                         in_data[305]
                    }),
            .out_data(lut_690_out)
        );

reg   lut_690_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_690_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_690_ff <= lut_690_out;
    end
end

assign out_data[690] = lut_690_ff;




// LUT : 691

wire lut_691_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101101000111111000010101011100011001001001001011111101011111),
            .DEVICE(DEVICE)
        )
    i_lut_691
        (
            .in_data({
                         in_data[40],
                         in_data[643],
                         in_data[107],
                         in_data[181],
                         in_data[551],
                         in_data[242]
                    }),
            .out_data(lut_691_out)
        );

reg   lut_691_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_691_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_691_ff <= lut_691_out;
    end
end

assign out_data[691] = lut_691_ff;




// LUT : 692

wire lut_692_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000111111000000101001011001001000111010000110010111101010010),
            .DEVICE(DEVICE)
        )
    i_lut_692
        (
            .in_data({
                         in_data[461],
                         in_data[626],
                         in_data[155],
                         in_data[3],
                         in_data[2],
                         in_data[59]
                    }),
            .out_data(lut_692_out)
        );

reg   lut_692_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_692_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_692_ff <= lut_692_out;
    end
end

assign out_data[692] = lut_692_ff;




// LUT : 693

wire lut_693_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111100000101001000011000100100001101011011011010111101010011),
            .DEVICE(DEVICE)
        )
    i_lut_693
        (
            .in_data({
                         in_data[400],
                         in_data[150],
                         in_data[153],
                         in_data[104],
                         in_data[624],
                         in_data[672]
                    }),
            .out_data(lut_693_out)
        );

reg   lut_693_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_693_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_693_ff <= lut_693_out;
    end
end

assign out_data[693] = lut_693_ff;




// LUT : 694

wire lut_694_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010011010110011101010111111001000000100110101101110101011110000),
            .DEVICE(DEVICE)
        )
    i_lut_694
        (
            .in_data({
                         in_data[439],
                         in_data[719],
                         in_data[648],
                         in_data[659],
                         in_data[186],
                         in_data[535]
                    }),
            .out_data(lut_694_out)
        );

reg   lut_694_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_694_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_694_ff <= lut_694_out;
    end
end

assign out_data[694] = lut_694_ff;




// LUT : 695

wire lut_695_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010001100110010011110011111100011100010010101011000100000000),
            .DEVICE(DEVICE)
        )
    i_lut_695
        (
            .in_data({
                         in_data[428],
                         in_data[753],
                         in_data[57],
                         in_data[238],
                         in_data[212],
                         in_data[601]
                    }),
            .out_data(lut_695_out)
        );

reg   lut_695_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_695_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_695_ff <= lut_695_out;
    end
end

assign out_data[695] = lut_695_ff;




// LUT : 696

wire lut_696_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110110010101110000000111001101111001110101101001100011111111111),
            .DEVICE(DEVICE)
        )
    i_lut_696
        (
            .in_data({
                         in_data[114],
                         in_data[389],
                         in_data[224],
                         in_data[654],
                         in_data[135],
                         in_data[276]
                    }),
            .out_data(lut_696_out)
        );

reg   lut_696_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_696_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_696_ff <= lut_696_out;
    end
end

assign out_data[696] = lut_696_ff;




// LUT : 697

wire lut_697_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010111111101100000100110110000100010010111100000100000100100001),
            .DEVICE(DEVICE)
        )
    i_lut_697
        (
            .in_data({
                         in_data[412],
                         in_data[425],
                         in_data[5],
                         in_data[71],
                         in_data[733],
                         in_data[120]
                    }),
            .out_data(lut_697_out)
        );

reg   lut_697_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_697_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_697_ff <= lut_697_out;
    end
end

assign out_data[697] = lut_697_ff;




// LUT : 698

wire lut_698_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001110110010100010010100010111100111001000100101110100000110101),
            .DEVICE(DEVICE)
        )
    i_lut_698
        (
            .in_data({
                         in_data[483],
                         in_data[721],
                         in_data[65],
                         in_data[113],
                         in_data[658],
                         in_data[162]
                    }),
            .out_data(lut_698_out)
        );

reg   lut_698_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_698_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_698_ff <= lut_698_out;
    end
end

assign out_data[698] = lut_698_ff;




// LUT : 699

wire lut_699_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001011000111100110011000001101011100101101110001101111110111101),
            .DEVICE(DEVICE)
        )
    i_lut_699
        (
            .in_data({
                         in_data[696],
                         in_data[645],
                         in_data[148],
                         in_data[142],
                         in_data[499],
                         in_data[364]
                    }),
            .out_data(lut_699_out)
        );

reg   lut_699_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_699_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_699_ff <= lut_699_out;
    end
end

assign out_data[699] = lut_699_ff;




// LUT : 700

wire lut_700_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111101100100000011011010010000011001000111000010010101110111101),
            .DEVICE(DEVICE)
        )
    i_lut_700
        (
            .in_data({
                         in_data[444],
                         in_data[702],
                         in_data[424],
                         in_data[669],
                         in_data[372],
                         in_data[174]
                    }),
            .out_data(lut_700_out)
        );

reg   lut_700_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_700_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_700_ff <= lut_700_out;
    end
end

assign out_data[700] = lut_700_ff;




// LUT : 701

wire lut_701_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100111011001111010101111101111010110011010111111011101101011110),
            .DEVICE(DEVICE)
        )
    i_lut_701
        (
            .in_data({
                         in_data[602],
                         in_data[415],
                         in_data[39],
                         in_data[628],
                         in_data[201],
                         in_data[68]
                    }),
            .out_data(lut_701_out)
        );

reg   lut_701_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_701_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_701_ff <= lut_701_out;
    end
end

assign out_data[701] = lut_701_ff;




// LUT : 702

wire lut_702_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010110010100011000111000011100101100001010011110001100101111),
            .DEVICE(DEVICE)
        )
    i_lut_702
        (
            .in_data({
                         in_data[296],
                         in_data[252],
                         in_data[320],
                         in_data[448],
                         in_data[95],
                         in_data[141]
                    }),
            .out_data(lut_702_out)
        );

reg   lut_702_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_702_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_702_ff <= lut_702_out;
    end
end

assign out_data[702] = lut_702_ff;




// LUT : 703

wire lut_703_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111111111100000111000001110010011110000),
            .DEVICE(DEVICE)
        )
    i_lut_703
        (
            .in_data({
                         in_data[525],
                         in_data[342],
                         in_data[341],
                         in_data[377],
                         in_data[687],
                         in_data[378]
                    }),
            .out_data(lut_703_out)
        );

reg   lut_703_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_703_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_703_ff <= lut_703_out;
    end
end

assign out_data[703] = lut_703_ff;




// LUT : 704

wire lut_704_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110001100000010110011001010011111111110111101111111111110100),
            .DEVICE(DEVICE)
        )
    i_lut_704
        (
            .in_data({
                         in_data[199],
                         in_data[442],
                         in_data[369],
                         in_data[291],
                         in_data[98],
                         in_data[128]
                    }),
            .out_data(lut_704_out)
        );

reg   lut_704_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_704_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_704_ff <= lut_704_out;
    end
end

assign out_data[704] = lut_704_ff;




// LUT : 705

wire lut_705_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111111011111110111010010101011111111010010100011000110101011),
            .DEVICE(DEVICE)
        )
    i_lut_705
        (
            .in_data({
                         in_data[72],
                         in_data[11],
                         in_data[339],
                         in_data[472],
                         in_data[180],
                         in_data[14]
                    }),
            .out_data(lut_705_out)
        );

reg   lut_705_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_705_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_705_ff <= lut_705_out;
    end
end

assign out_data[705] = lut_705_ff;




// LUT : 706

wire lut_706_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111101100111011001001101111111011101001001110000100011101010),
            .DEVICE(DEVICE)
        )
    i_lut_706
        (
            .in_data({
                         in_data[457],
                         in_data[330],
                         in_data[594],
                         in_data[383],
                         in_data[430],
                         in_data[23]
                    }),
            .out_data(lut_706_out)
        );

reg   lut_706_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_706_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_706_ff <= lut_706_out;
    end
end

assign out_data[706] = lut_706_ff;




// LUT : 707

wire lut_707_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001011111010011010111111101001110010000100000000011111111011),
            .DEVICE(DEVICE)
        )
    i_lut_707
        (
            .in_data({
                         in_data[152],
                         in_data[189],
                         in_data[423],
                         in_data[92],
                         in_data[527],
                         in_data[268]
                    }),
            .out_data(lut_707_out)
        );

reg   lut_707_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_707_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_707_ff <= lut_707_out;
    end
end

assign out_data[707] = lut_707_ff;




// LUT : 708

wire lut_708_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001111010011000100001001010101101000000111011110010011010100101),
            .DEVICE(DEVICE)
        )
    i_lut_708
        (
            .in_data({
                         in_data[15],
                         in_data[636],
                         in_data[599],
                         in_data[519],
                         in_data[286],
                         in_data[367]
                    }),
            .out_data(lut_708_out)
        );

reg   lut_708_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_708_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_708_ff <= lut_708_out;
    end
end

assign out_data[708] = lut_708_ff;




// LUT : 709

wire lut_709_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101111000001101110001110011110000100011000001100110011010110),
            .DEVICE(DEVICE)
        )
    i_lut_709
        (
            .in_data({
                         in_data[43],
                         in_data[119],
                         in_data[49],
                         in_data[157],
                         in_data[664],
                         in_data[54]
                    }),
            .out_data(lut_709_out)
        );

reg   lut_709_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_709_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_709_ff <= lut_709_out;
    end
end

assign out_data[709] = lut_709_ff;




// LUT : 710

wire lut_710_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000001011001111010000010101000000100001100000000000010000010),
            .DEVICE(DEVICE)
        )
    i_lut_710
        (
            .in_data({
                         in_data[132],
                         in_data[610],
                         in_data[282],
                         in_data[311],
                         in_data[711],
                         in_data[635]
                    }),
            .out_data(lut_710_out)
        );

reg   lut_710_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_710_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_710_ff <= lut_710_out;
    end
end

assign out_data[710] = lut_710_ff;




// LUT : 711

wire lut_711_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111100001111101000100111100011111011001101100010001100000010001),
            .DEVICE(DEVICE)
        )
    i_lut_711
        (
            .in_data({
                         in_data[30],
                         in_data[158],
                         in_data[600],
                         in_data[522],
                         in_data[354],
                         in_data[112]
                    }),
            .out_data(lut_711_out)
        );

reg   lut_711_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_711_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_711_ff <= lut_711_out;
    end
end

assign out_data[711] = lut_711_ff;




// LUT : 712

wire lut_712_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000010110001011000000111110001000101001011010110000100000001),
            .DEVICE(DEVICE)
        )
    i_lut_712
        (
            .in_data({
                         in_data[47],
                         in_data[651],
                         in_data[403],
                         in_data[587],
                         in_data[134],
                         in_data[164]
                    }),
            .out_data(lut_712_out)
        );

reg   lut_712_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_712_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_712_ff <= lut_712_out;
    end
end

assign out_data[712] = lut_712_ff;




// LUT : 713

wire lut_713_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100000100010110011001100100011001100101010101100111111101111),
            .DEVICE(DEVICE)
        )
    i_lut_713
        (
            .in_data({
                         in_data[481],
                         in_data[580],
                         in_data[453],
                         in_data[577],
                         in_data[414],
                         in_data[486]
                    }),
            .out_data(lut_713_out)
        );

reg   lut_713_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_713_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_713_ff <= lut_713_out;
    end
end

assign out_data[713] = lut_713_ff;




// LUT : 714

wire lut_714_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010100010111010111010111110111000110011111110011000001110100),
            .DEVICE(DEVICE)
        )
    i_lut_714
        (
            .in_data({
                         in_data[353],
                         in_data[730],
                         in_data[598],
                         in_data[409],
                         in_data[355],
                         in_data[241]
                    }),
            .out_data(lut_714_out)
        );

reg   lut_714_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_714_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_714_ff <= lut_714_out;
    end
end

assign out_data[714] = lut_714_ff;




// LUT : 715

wire lut_715_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010010000000000111110111000000011011010000011001100101101001101),
            .DEVICE(DEVICE)
        )
    i_lut_715
        (
            .in_data({
                         in_data[185],
                         in_data[489],
                         in_data[85],
                         in_data[243],
                         in_data[410],
                         in_data[387]
                    }),
            .out_data(lut_715_out)
        );

reg   lut_715_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_715_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_715_ff <= lut_715_out;
    end
end

assign out_data[715] = lut_715_ff;




// LUT : 716

wire lut_716_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010011101111001000010110010010110001111011110101000000000100100),
            .DEVICE(DEVICE)
        )
    i_lut_716
        (
            .in_data({
                         in_data[284],
                         in_data[255],
                         in_data[402],
                         in_data[737],
                         in_data[365],
                         in_data[106]
                    }),
            .out_data(lut_716_out)
        );

reg   lut_716_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_716_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_716_ff <= lut_716_out;
    end
end

assign out_data[716] = lut_716_ff;




// LUT : 717

wire lut_717_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101001111101111001000011000011100100101111010110100000101100011),
            .DEVICE(DEVICE)
        )
    i_lut_717
        (
            .in_data({
                         in_data[653],
                         in_data[739],
                         in_data[515],
                         in_data[223],
                         in_data[556],
                         in_data[455]
                    }),
            .out_data(lut_717_out)
        );

reg   lut_717_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_717_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_717_ff <= lut_717_out;
    end
end

assign out_data[717] = lut_717_ff;




// LUT : 718

wire lut_718_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000101000110001010111111101100110000001000111111100000111011),
            .DEVICE(DEVICE)
        )
    i_lut_718
        (
            .in_data({
                         in_data[101],
                         in_data[662],
                         in_data[208],
                         in_data[244],
                         in_data[504],
                         in_data[668]
                    }),
            .out_data(lut_718_out)
        );

reg   lut_718_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_718_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_718_ff <= lut_718_out;
    end
end

assign out_data[718] = lut_718_ff;




// LUT : 719

wire lut_719_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100001010001100010001001000100000100000011000001010101011001),
            .DEVICE(DEVICE)
        )
    i_lut_719
        (
            .in_data({
                         in_data[682],
                         in_data[688],
                         in_data[540],
                         in_data[583],
                         in_data[16],
                         in_data[302]
                    }),
            .out_data(lut_719_out)
        );

reg   lut_719_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_719_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_719_ff <= lut_719_out;
    end
end

assign out_data[719] = lut_719_ff;




// LUT : 720

wire lut_720_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010101110010001011010001010011001010111001001111100101011001),
            .DEVICE(DEVICE)
        )
    i_lut_720
        (
            .in_data({
                         in_data[29],
                         in_data[530],
                         in_data[652],
                         in_data[136],
                         in_data[206],
                         in_data[22]
                    }),
            .out_data(lut_720_out)
        );

reg   lut_720_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_720_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_720_ff <= lut_720_out;
    end
end

assign out_data[720] = lut_720_ff;




// LUT : 721

wire lut_721_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100110001011011000001100110001000110000101001110010101100100),
            .DEVICE(DEVICE)
        )
    i_lut_721
        (
            .in_data({
                         in_data[12],
                         in_data[171],
                         in_data[440],
                         in_data[281],
                         in_data[357],
                         in_data[720]
                    }),
            .out_data(lut_721_out)
        );

reg   lut_721_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_721_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_721_ff <= lut_721_out;
    end
end

assign out_data[721] = lut_721_ff;




// LUT : 722

wire lut_722_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111111110011010111001001000101110011001101000011010000101100),
            .DEVICE(DEVICE)
        )
    i_lut_722
        (
            .in_data({
                         in_data[118],
                         in_data[126],
                         in_data[325],
                         in_data[173],
                         in_data[366],
                         in_data[468]
                    }),
            .out_data(lut_722_out)
        );

reg   lut_722_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_722_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_722_ff <= lut_722_out;
    end
end

assign out_data[722] = lut_722_ff;




// LUT : 723

wire lut_723_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010010100101011011000001000111011111001001000001111000010001),
            .DEVICE(DEVICE)
        )
    i_lut_723
        (
            .in_data({
                         in_data[488],
                         in_data[10],
                         in_data[673],
                         in_data[347],
                         in_data[231],
                         in_data[257]
                    }),
            .out_data(lut_723_out)
        );

reg   lut_723_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_723_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_723_ff <= lut_723_out;
    end
end

assign out_data[723] = lut_723_ff;




// LUT : 724

wire lut_724_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110110101110011111110101011011101001100101110111111000001101100),
            .DEVICE(DEVICE)
        )
    i_lut_724
        (
            .in_data({
                         in_data[557],
                         in_data[445],
                         in_data[219],
                         in_data[686],
                         in_data[394],
                         in_data[348]
                    }),
            .out_data(lut_724_out)
        );

reg   lut_724_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_724_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_724_ff <= lut_724_out;
    end
end

assign out_data[724] = lut_724_ff;




// LUT : 725

wire lut_725_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101000110011101000000011000010111111111110111111000011110000),
            .DEVICE(DEVICE)
        )
    i_lut_725
        (
            .in_data({
                         in_data[319],
                         in_data[581],
                         in_data[573],
                         in_data[151],
                         in_data[316],
                         in_data[517]
                    }),
            .out_data(lut_725_out)
        );

reg   lut_725_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_725_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_725_ff <= lut_725_out;
    end
end

assign out_data[725] = lut_725_ff;




// LUT : 726

wire lut_726_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100011000011100000110100100010100000011000111111011011001100),
            .DEVICE(DEVICE)
        )
    i_lut_726
        (
            .in_data({
                         in_data[735],
                         in_data[478],
                         in_data[533],
                         in_data[299],
                         in_data[83],
                         in_data[411]
                    }),
            .out_data(lut_726_out)
        );

reg   lut_726_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_726_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_726_ff <= lut_726_out;
    end
end

assign out_data[726] = lut_726_ff;




// LUT : 727

wire lut_727_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110101111111111101011011110111110011101001000011111101100100),
            .DEVICE(DEVICE)
        )
    i_lut_727
        (
            .in_data({
                         in_data[338],
                         in_data[379],
                         in_data[266],
                         in_data[500],
                         in_data[310],
                         in_data[358]
                    }),
            .out_data(lut_727_out)
        );

reg   lut_727_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_727_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_727_ff <= lut_727_out;
    end
end

assign out_data[727] = lut_727_ff;




// LUT : 728

wire lut_728_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111010100101011101001110000010100000110001111011010000101000),
            .DEVICE(DEVICE)
        )
    i_lut_728
        (
            .in_data({
                         in_data[431],
                         in_data[529],
                         in_data[218],
                         in_data[619],
                         in_data[99],
                         in_data[35]
                    }),
            .out_data(lut_728_out)
        );

reg   lut_728_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_728_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_728_ff <= lut_728_out;
    end
end

assign out_data[728] = lut_728_ff;




// LUT : 729

wire lut_729_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011011111111101111101011011111111110101011110011110100000000),
            .DEVICE(DEVICE)
        )
    i_lut_729
        (
            .in_data({
                         in_data[490],
                         in_data[109],
                         in_data[38],
                         in_data[396],
                         in_data[544],
                         in_data[482]
                    }),
            .out_data(lut_729_out)
        );

reg   lut_729_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_729_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_729_ff <= lut_729_out;
    end
end

assign out_data[729] = lut_729_ff;




// LUT : 730

wire lut_730_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010100000101101111111101001011101111111111011010001011011011),
            .DEVICE(DEVICE)
        )
    i_lut_730
        (
            .in_data({
                         in_data[392],
                         in_data[87],
                         in_data[596],
                         in_data[712],
                         in_data[270],
                         in_data[703]
                    }),
            .out_data(lut_730_out)
        );

reg   lut_730_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_730_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_730_ff <= lut_730_out;
    end
end

assign out_data[730] = lut_730_ff;




// LUT : 731

wire lut_731_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110010101010100111101000101101101000100010010000011001000101),
            .DEVICE(DEVICE)
        )
    i_lut_731
        (
            .in_data({
                         in_data[24],
                         in_data[752],
                         in_data[247],
                         in_data[476],
                         in_data[505],
                         in_data[88]
                    }),
            .out_data(lut_731_out)
        );

reg   lut_731_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_731_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_731_ff <= lut_731_out;
    end
end

assign out_data[731] = lut_731_ff;




// LUT : 732

wire lut_732_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001011000110101011110100110110100000011000100000101001000100),
            .DEVICE(DEVICE)
        )
    i_lut_732
        (
            .in_data({
                         in_data[216],
                         in_data[331],
                         in_data[234],
                         in_data[595],
                         in_data[260],
                         in_data[675]
                    }),
            .out_data(lut_732_out)
        );

reg   lut_732_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_732_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_732_ff <= lut_732_out;
    end
end

assign out_data[732] = lut_732_ff;




// LUT : 733

wire lut_733_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000001000101101100001000100000000000000001010101001111001101),
            .DEVICE(DEVICE)
        )
    i_lut_733
        (
            .in_data({
                         in_data[484],
                         in_data[516],
                         in_data[563],
                         in_data[612],
                         in_data[441],
                         in_data[541]
                    }),
            .out_data(lut_733_out)
        );

reg   lut_733_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_733_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_733_ff <= lut_733_out;
    end
end

assign out_data[733] = lut_733_ff;




// LUT : 734

wire lut_734_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110010101000000100001110100000010001011100011000000100001001),
            .DEVICE(DEVICE)
        )
    i_lut_734
        (
            .in_data({
                         in_data[692],
                         in_data[497],
                         in_data[460],
                         in_data[363],
                         in_data[683],
                         in_data[724]
                    }),
            .out_data(lut_734_out)
        );

reg   lut_734_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_734_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_734_ff <= lut_734_out;
    end
end

assign out_data[734] = lut_734_ff;




// LUT : 735

wire lut_735_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111001010010001110100101111100111010111110100111010000110100),
            .DEVICE(DEVICE)
        )
    i_lut_735
        (
            .in_data({
                         in_data[552],
                         in_data[329],
                         in_data[124],
                         in_data[121],
                         in_data[644],
                         in_data[432]
                    }),
            .out_data(lut_735_out)
        );

reg   lut_735_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_735_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_735_ff <= lut_735_out;
    end
end

assign out_data[735] = lut_735_ff;




// LUT : 736

wire lut_736_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001101011111000110000110010111011110111101000101110111111110),
            .DEVICE(DEVICE)
        )
    i_lut_736
        (
            .in_data({
                         in_data[306],
                         in_data[707],
                         in_data[160],
                         in_data[701],
                         in_data[605],
                         in_data[125]
                    }),
            .out_data(lut_736_out)
        );

reg   lut_736_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_736_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_736_ff <= lut_736_out;
    end
end

assign out_data[736] = lut_736_ff;




// LUT : 737

wire lut_737_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000100101000000000001000001000000000100010000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_737
        (
            .in_data({
                         in_data[249],
                         in_data[561],
                         in_data[492],
                         in_data[401],
                         in_data[382],
                         in_data[67]
                    }),
            .out_data(lut_737_out)
        );

reg   lut_737_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_737_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_737_ff <= lut_737_out;
    end
end

assign out_data[737] = lut_737_ff;




// LUT : 738

wire lut_738_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010010110001101001001000100110000010111101111010110000001111111),
            .DEVICE(DEVICE)
        )
    i_lut_738
        (
            .in_data({
                         in_data[381],
                         in_data[333],
                         in_data[388],
                         in_data[778],
                         in_data[568],
                         in_data[137]
                    }),
            .out_data(lut_738_out)
        );

reg   lut_738_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_738_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_738_ff <= lut_738_out;
    end
end

assign out_data[738] = lut_738_ff;




// LUT : 739

wire lut_739_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000101111010000100001000100011011101010100001101100101101001),
            .DEVICE(DEVICE)
        )
    i_lut_739
        (
            .in_data({
                         in_data[463],
                         in_data[41],
                         in_data[293],
                         in_data[117],
                         in_data[501],
                         in_data[507]
                    }),
            .out_data(lut_739_out)
        );

reg   lut_739_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_739_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_739_ff <= lut_739_out;
    end
end

assign out_data[739] = lut_739_ff;




// LUT : 740

wire lut_740_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001101110111111110111111110101000011110111100111101110100111110),
            .DEVICE(DEVICE)
        )
    i_lut_740
        (
            .in_data({
                         in_data[465],
                         in_data[309],
                         in_data[89],
                         in_data[633],
                         in_data[335],
                         in_data[263]
                    }),
            .out_data(lut_740_out)
        );

reg   lut_740_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_740_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_740_ff <= lut_740_out;
    end
end

assign out_data[740] = lut_740_ff;




// LUT : 741

wire lut_741_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101010110100111111010110110111110100111011010111011100001110),
            .DEVICE(DEVICE)
        )
    i_lut_741
        (
            .in_data({
                         in_data[225],
                         in_data[248],
                         in_data[205],
                         in_data[362],
                         in_data[649],
                         in_data[479]
                    }),
            .out_data(lut_741_out)
        );

reg   lut_741_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_741_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_741_ff <= lut_741_out;
    end
end

assign out_data[741] = lut_741_ff;




// LUT : 742

wire lut_742_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000010110100000000011100100110011010100000000110110011001101),
            .DEVICE(DEVICE)
        )
    i_lut_742
        (
            .in_data({
                         in_data[655],
                         in_data[582],
                         in_data[717],
                         in_data[69],
                         in_data[700],
                         in_data[221]
                    }),
            .out_data(lut_742_out)
        );

reg   lut_742_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_742_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_742_ff <= lut_742_out;
    end
end

assign out_data[742] = lut_742_ff;




// LUT : 743

wire lut_743_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110101001110010110001100010000000111000001000100110000010011),
            .DEVICE(DEVICE)
        )
    i_lut_743
        (
            .in_data({
                         in_data[386],
                         in_data[32],
                         in_data[45],
                         in_data[93],
                         in_data[742],
                         in_data[262]
                    }),
            .out_data(lut_743_out)
        );

reg   lut_743_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_743_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_743_ff <= lut_743_out;
    end
end

assign out_data[743] = lut_743_ff;




// LUT : 744

wire lut_744_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100111110010000010001110011110111011101010011110011000011101101),
            .DEVICE(DEVICE)
        )
    i_lut_744
        (
            .in_data({
                         in_data[307],
                         in_data[96],
                         in_data[323],
                         in_data[60],
                         in_data[547],
                         in_data[443]
                    }),
            .out_data(lut_744_out)
        );

reg   lut_744_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_744_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_744_ff <= lut_744_out;
    end
end

assign out_data[744] = lut_744_ff;




// LUT : 745

wire lut_745_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110000001101000010100100000111010011001110011111111110111000011),
            .DEVICE(DEVICE)
        )
    i_lut_745
        (
            .in_data({
                         in_data[741],
                         in_data[511],
                         in_data[308],
                         in_data[73],
                         in_data[780],
                         in_data[565]
                    }),
            .out_data(lut_745_out)
        );

reg   lut_745_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_745_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_745_ff <= lut_745_out;
    end
end

assign out_data[745] = lut_745_ff;




// LUT : 746

wire lut_746_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100101010111011011011111110110011101101101011101110011111111),
            .DEVICE(DEVICE)
        )
    i_lut_746
        (
            .in_data({
                         in_data[546],
                         in_data[487],
                         in_data[614],
                         in_data[251],
                         in_data[192],
                         in_data[592]
                    }),
            .out_data(lut_746_out)
        );

reg   lut_746_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_746_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_746_ff <= lut_746_out;
    end
end

assign out_data[746] = lut_746_ff;




// LUT : 747

wire lut_747_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100010010100100001111100100000111100001000011000110110110000101),
            .DEVICE(DEVICE)
        )
    i_lut_747
        (
            .in_data({
                         in_data[661],
                         in_data[90],
                         in_data[390],
                         in_data[708],
                         in_data[666],
                         in_data[261]
                    }),
            .out_data(lut_747_out)
        );

reg   lut_747_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_747_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_747_ff <= lut_747_out;
    end
end

assign out_data[747] = lut_747_ff;




// LUT : 748

wire lut_748_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100111100101011011110110110111100111110100111101100110001111100),
            .DEVICE(DEVICE)
        )
    i_lut_748
        (
            .in_data({
                         in_data[763],
                         in_data[710],
                         in_data[520],
                         in_data[18],
                         in_data[480],
                         in_data[606]
                    }),
            .out_data(lut_748_out)
        );

reg   lut_748_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_748_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_748_ff <= lut_748_out;
    end
end

assign out_data[748] = lut_748_ff;




// LUT : 749

wire lut_749_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010110011001100101011011110101100101011000000000010101100000),
            .DEVICE(DEVICE)
        )
    i_lut_749
        (
            .in_data({
                         in_data[715],
                         in_data[376],
                         in_data[631],
                         in_data[781],
                         in_data[328],
                         in_data[684]
                    }),
            .out_data(lut_749_out)
        );

reg   lut_749_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_749_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_749_ff <= lut_749_out;
    end
end

assign out_data[749] = lut_749_ff;




// LUT : 750

wire lut_750_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111010110111011010100001100101101000001101101100000011101110),
            .DEVICE(DEVICE)
        )
    i_lut_750
        (
            .in_data({
                         in_data[538],
                         in_data[622],
                         in_data[417],
                         in_data[604],
                         in_data[757],
                         in_data[618]
                    }),
            .out_data(lut_750_out)
        );

reg   lut_750_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_750_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_750_ff <= lut_750_out;
    end
end

assign out_data[750] = lut_750_ff;




// LUT : 751

wire lut_751_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011110100111011101110011111111100100010001110101101010011001100),
            .DEVICE(DEVICE)
        )
    i_lut_751
        (
            .in_data({
                         in_data[368],
                         in_data[214],
                         in_data[217],
                         in_data[466],
                         in_data[671],
                         in_data[264]
                    }),
            .out_data(lut_751_out)
        );

reg   lut_751_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_751_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_751_ff <= lut_751_out;
    end
end

assign out_data[751] = lut_751_ff;




// LUT : 752

wire lut_752_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100011110100111011101010001101010011011000110001010110000110),
            .DEVICE(DEVICE)
        )
    i_lut_752
        (
            .in_data({
                         in_data[782],
                         in_data[759],
                         in_data[681],
                         in_data[345],
                         in_data[508],
                         in_data[391]
                    }),
            .out_data(lut_752_out)
        );

reg   lut_752_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_752_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_752_ff <= lut_752_out;
    end
end

assign out_data[752] = lut_752_ff;




// LUT : 753

wire lut_753_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010011001100010100001110101010001101100011101100011000101001),
            .DEVICE(DEVICE)
        )
    i_lut_753
        (
            .in_data({
                         in_data[190],
                         in_data[385],
                         in_data[200],
                         in_data[413],
                         in_data[760],
                         in_data[526]
                    }),
            .out_data(lut_753_out)
        );

reg   lut_753_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_753_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_753_ff <= lut_753_out;
    end
end

assign out_data[753] = lut_753_ff;




// LUT : 754

wire lut_754_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000100001111001110110100111000100100111011011001001111110110),
            .DEVICE(DEVICE)
        )
    i_lut_754
        (
            .in_data({
                         in_data[240],
                         in_data[734],
                         in_data[165],
                         in_data[227],
                         in_data[764],
                         in_data[694]
                    }),
            .out_data(lut_754_out)
        );

reg   lut_754_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_754_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_754_ff <= lut_754_out;
    end
end

assign out_data[754] = lut_754_ff;




// LUT : 755

wire lut_755_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111110010100110111001010010101111001100110101000100001100010011),
            .DEVICE(DEVICE)
        )
    i_lut_755
        (
            .in_data({
                         in_data[56],
                         in_data[674],
                         in_data[532],
                         in_data[471],
                         in_data[75],
                         in_data[374]
                    }),
            .out_data(lut_755_out)
        );

reg   lut_755_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_755_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_755_ff <= lut_755_out;
    end
end

assign out_data[755] = lut_755_ff;




// LUT : 756

wire lut_756_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001111110101110100110001000101001100100111000011011101110000),
            .DEVICE(DEVICE)
        )
    i_lut_756
        (
            .in_data({
                         in_data[337],
                         in_data[464],
                         in_data[743],
                         in_data[313],
                         in_data[726],
                         in_data[294]
                    }),
            .out_data(lut_756_out)
        );

reg   lut_756_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_756_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_756_ff <= lut_756_out;
    end
end

assign out_data[756] = lut_756_ff;




// LUT : 757

wire lut_757_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001011010100000000111111100000001001111011111001110011100001),
            .DEVICE(DEVICE)
        )
    i_lut_757
        (
            .in_data({
                         in_data[779],
                         in_data[722],
                         in_data[61],
                         in_data[7],
                         in_data[593],
                         in_data[230]
                    }),
            .out_data(lut_757_out)
        );

reg   lut_757_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_757_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_757_ff <= lut_757_out;
    end
end

assign out_data[757] = lut_757_ff;




// LUT : 758

wire lut_758_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000011100111111001000111000011100010000010000101001110010000),
            .DEVICE(DEVICE)
        )
    i_lut_758
        (
            .in_data({
                         in_data[680],
                         in_data[370],
                         in_data[84],
                         in_data[698],
                         in_data[616],
                         in_data[167]
                    }),
            .out_data(lut_758_out)
        );

reg   lut_758_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_758_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_758_ff <= lut_758_out;
    end
end

assign out_data[758] = lut_758_ff;




// LUT : 759

wire lut_759_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100101100100101000001001101100000100000100001000010000010001),
            .DEVICE(DEVICE)
        )
    i_lut_759
        (
            .in_data({
                         in_data[736],
                         in_data[177],
                         in_data[116],
                         in_data[322],
                         in_data[677],
                         in_data[657]
                    }),
            .out_data(lut_759_out)
        );

reg   lut_759_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_759_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_759_ff <= lut_759_out;
    end
end

assign out_data[759] = lut_759_ff;




// LUT : 760

wire lut_760_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001100100000110111110010010111001001101010001001010011101100010),
            .DEVICE(DEVICE)
        )
    i_lut_760
        (
            .in_data({
                         in_data[650],
                         in_data[274],
                         in_data[349],
                         in_data[318],
                         in_data[758],
                         in_data[166]
                    }),
            .out_data(lut_760_out)
        );

reg   lut_760_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_760_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_760_ff <= lut_760_out;
    end
end

assign out_data[760] = lut_760_ff;




// LUT : 761

wire lut_761_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111111111111011001101010000010000000110100001000101100000011),
            .DEVICE(DEVICE)
        )
    i_lut_761
        (
            .in_data({
                         in_data[62],
                         in_data[783],
                         in_data[549],
                         in_data[127],
                         in_data[474],
                         in_data[705]
                    }),
            .out_data(lut_761_out)
        );

reg   lut_761_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_761_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_761_ff <= lut_761_out;
    end
end

assign out_data[761] = lut_761_ff;




// LUT : 762

wire lut_762_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101100101110110110010011111011100000010111111111000000000111100),
            .DEVICE(DEVICE)
        )
    i_lut_762
        (
            .in_data({
                         in_data[713],
                         in_data[718],
                         in_data[6],
                         in_data[344],
                         in_data[395],
                         in_data[553]
                    }),
            .out_data(lut_762_out)
        );

reg   lut_762_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_762_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_762_ff <= lut_762_out;
    end
end

assign out_data[762] = lut_762_ff;




// LUT : 763

wire lut_763_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100110111011111111111011111011010111111101111111111111101100),
            .DEVICE(DEVICE)
        )
    i_lut_763
        (
            .in_data({
                         in_data[371],
                         in_data[91],
                         in_data[427],
                         in_data[100],
                         in_data[191],
                         in_data[433]
                    }),
            .out_data(lut_763_out)
        );

reg   lut_763_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_763_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_763_ff <= lut_763_out;
    end
end

assign out_data[763] = lut_763_ff;




// LUT : 764

wire lut_764_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100011001100010000100111111111111000101011000101010101101000),
            .DEVICE(DEVICE)
        )
    i_lut_764
        (
            .in_data({
                         in_data[278],
                         in_data[404],
                         in_data[523],
                         in_data[531],
                         in_data[28],
                         in_data[146]
                    }),
            .out_data(lut_764_out)
        );

reg   lut_764_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_764_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_764_ff <= lut_764_out;
    end
end

assign out_data[764] = lut_764_ff;




// LUT : 765

wire lut_765_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101000101011011010101100000110110111011011001000011000010101),
            .DEVICE(DEVICE)
        )
    i_lut_765
        (
            .in_data({
                         in_data[745],
                         in_data[129],
                         in_data[744],
                         in_data[235],
                         in_data[560],
                         in_data[559]
                    }),
            .out_data(lut_765_out)
        );

reg   lut_765_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_765_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_765_ff <= lut_765_out;
    end
end

assign out_data[765] = lut_765_ff;




// LUT : 766

wire lut_766_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001001000011000011101101100000001000100000010001011111000100001),
            .DEVICE(DEVICE)
        )
    i_lut_766
        (
            .in_data({
                         in_data[277],
                         in_data[534],
                         in_data[725],
                         in_data[178],
                         in_data[193],
                         in_data[586]
                    }),
            .out_data(lut_766_out)
        );

reg   lut_766_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_766_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_766_ff <= lut_766_out;
    end
end

assign out_data[766] = lut_766_ff;




// LUT : 767

wire lut_767_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110000000110110000001101001011001111001100011110011011011001),
            .DEVICE(DEVICE)
        )
    i_lut_767
        (
            .in_data({
                         in_data[754],
                         in_data[312],
                         in_data[48],
                         in_data[749],
                         in_data[194],
                         in_data[420]
                    }),
            .out_data(lut_767_out)
        );

reg   lut_767_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_767_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_767_ff <= lut_767_out;
    end
end

assign out_data[767] = lut_767_ff;




// LUT : 768

wire lut_768_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100111110010010111010000011111100011101000101111101010101110),
            .DEVICE(DEVICE)
        )
    i_lut_768
        (
            .in_data({
                         in_data[222],
                         in_data[279],
                         in_data[34],
                         in_data[435],
                         in_data[285],
                         in_data[131]
                    }),
            .out_data(lut_768_out)
        );

reg   lut_768_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_768_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_768_ff <= lut_768_out;
    end
end

assign out_data[768] = lut_768_ff;




// LUT : 769

wire lut_769_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111001000010001110100010100100011111001000001000001001110111),
            .DEVICE(DEVICE)
        )
    i_lut_769
        (
            .in_data({
                         in_data[336],
                         in_data[408],
                         in_data[55],
                         in_data[639],
                         in_data[350],
                         in_data[591]
                    }),
            .out_data(lut_769_out)
        );

reg   lut_769_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_769_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_769_ff <= lut_769_out;
    end
end

assign out_data[769] = lut_769_ff;




// LUT : 770

wire lut_770_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001111001010010011101110111010010110010011100000101001011010000),
            .DEVICE(DEVICE)
        )
    i_lut_770
        (
            .in_data({
                         in_data[346],
                         in_data[184],
                         in_data[558],
                         in_data[714],
                         in_data[297],
                         in_data[321]
                    }),
            .out_data(lut_770_out)
        );

reg   lut_770_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_770_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_770_ff <= lut_770_out;
    end
end

assign out_data[770] = lut_770_ff;




// LUT : 771

wire lut_771_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111101110011110011111010000010000010000101001011101010100100),
            .DEVICE(DEVICE)
        )
    i_lut_771
        (
            .in_data({
                         in_data[66],
                         in_data[81],
                         in_data[25],
                         in_data[416],
                         in_data[607],
                         in_data[280]
                    }),
            .out_data(lut_771_out)
        );

reg   lut_771_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_771_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_771_ff <= lut_771_out;
    end
end

assign out_data[771] = lut_771_ff;




// LUT : 772

wire lut_772_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010000101110010100000101101101000101011000010010010001010001),
            .DEVICE(DEVICE)
        )
    i_lut_772
        (
            .in_data({
                         in_data[245],
                         in_data[197],
                         in_data[304],
                         in_data[421],
                         in_data[762],
                         in_data[103]
                    }),
            .out_data(lut_772_out)
        );

reg   lut_772_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_772_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_772_ff <= lut_772_out;
    end
end

assign out_data[772] = lut_772_ff;




// LUT : 773

wire lut_773_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110110101010111010111111100111101101110010111110010111111011010),
            .DEVICE(DEVICE)
        )
    i_lut_773
        (
            .in_data({
                         in_data[536],
                         in_data[78],
                         in_data[665],
                         in_data[86],
                         in_data[288],
                         in_data[498]
                    }),
            .out_data(lut_773_out)
        );

reg   lut_773_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_773_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_773_ff <= lut_773_out;
    end
end

assign out_data[773] = lut_773_ff;




// LUT : 774

wire lut_774_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010010011101101010101110111101100001000000000000000000001100),
            .DEVICE(DEVICE)
        )
    i_lut_774
        (
            .in_data({
                         in_data[429],
                         in_data[678],
                         in_data[272],
                         in_data[298],
                         in_data[237],
                         in_data[290]
                    }),
            .out_data(lut_774_out)
        );

reg   lut_774_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_774_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_774_ff <= lut_774_out;
    end
end

assign out_data[774] = lut_774_ff;




// LUT : 775

wire lut_775_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111011110111100010000010001001100110110100001100111011010100),
            .DEVICE(DEVICE)
        )
    i_lut_775
        (
            .in_data({
                         in_data[510],
                         in_data[210],
                         in_data[777],
                         in_data[172],
                         in_data[198],
                         in_data[621]
                    }),
            .out_data(lut_775_out)
        );

reg   lut_775_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_775_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_775_ff <= lut_775_out;
    end
end

assign out_data[775] = lut_775_ff;




// LUT : 776

wire lut_776_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011010111100101010111011100111111101101001111111001101001010000),
            .DEVICE(DEVICE)
        )
    i_lut_776
        (
            .in_data({
                         in_data[447],
                         in_data[446],
                         in_data[470],
                         in_data[765],
                         in_data[373],
                         in_data[195]
                    }),
            .out_data(lut_776_out)
        );

reg   lut_776_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_776_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_776_ff <= lut_776_out;
    end
end

assign out_data[776] = lut_776_ff;




// LUT : 777

wire lut_777_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111111001101111111111111111111010000010000000011011111111011),
            .DEVICE(DEVICE)
        )
    i_lut_777
        (
            .in_data({
                         in_data[188],
                         in_data[295],
                         in_data[693],
                         in_data[467],
                         in_data[163],
                         in_data[690]
                    }),
            .out_data(lut_777_out)
        );

reg   lut_777_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_777_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_777_ff <= lut_777_out;
    end
end

assign out_data[777] = lut_777_ff;




// LUT : 778

wire lut_778_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011101111010110010011111010101011110011010000001010111001011100),
            .DEVICE(DEVICE)
        )
    i_lut_778
        (
            .in_data({
                         in_data[1],
                         in_data[327],
                         in_data[751],
                         in_data[130],
                         in_data[554],
                         in_data[283]
                    }),
            .out_data(lut_778_out)
        );

reg   lut_778_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_778_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_778_ff <= lut_778_out;
    end
end

assign out_data[778] = lut_778_ff;




// LUT : 779

wire lut_779_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100010010010111100000001100100011011100110000001000100001001001),
            .DEVICE(DEVICE)
        )
    i_lut_779
        (
            .in_data({
                         in_data[449],
                         in_data[496],
                         in_data[454],
                         in_data[584],
                         in_data[589],
                         in_data[585]
                    }),
            .out_data(lut_779_out)
        );

reg   lut_779_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_779_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_779_ff <= lut_779_out;
    end
end

assign out_data[779] = lut_779_ff;




// LUT : 780

wire lut_780_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001110111001011110011110101001010111100100011101010111111010),
            .DEVICE(DEVICE)
        )
    i_lut_780
        (
            .in_data({
                         in_data[509],
                         in_data[551],
                         in_data[361],
                         in_data[571],
                         in_data[300],
                         in_data[620]
                    }),
            .out_data(lut_780_out)
        );

reg   lut_780_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_780_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_780_ff <= lut_780_out;
    end
end

assign out_data[780] = lut_780_ff;




// LUT : 781

wire lut_781_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001001111110001101110110111110000010000111111011010111111111),
            .DEVICE(DEVICE)
        )
    i_lut_781
        (
            .in_data({
                         in_data[756],
                         in_data[697],
                         in_data[449],
                         in_data[397],
                         in_data[170],
                         in_data[33]
                    }),
            .out_data(lut_781_out)
        );

reg   lut_781_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_781_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_781_ff <= lut_781_out;
    end
end

assign out_data[781] = lut_781_ff;




// LUT : 782

wire lut_782_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000000100100010000001010011011010100101000000011001101011101),
            .DEVICE(DEVICE)
        )
    i_lut_782
        (
            .in_data({
                         in_data[485],
                         in_data[194],
                         in_data[184],
                         in_data[562],
                         in_data[779],
                         in_data[614]
                    }),
            .out_data(lut_782_out)
        );

reg   lut_782_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_782_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_782_ff <= lut_782_out;
    end
end

assign out_data[782] = lut_782_ff;




// LUT : 783

wire lut_783_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000100010111000000011011101110010100110010001011010000000000),
            .DEVICE(DEVICE)
        )
    i_lut_783
        (
            .in_data({
                         in_data[352],
                         in_data[427],
                         in_data[111],
                         in_data[603],
                         in_data[52],
                         in_data[215]
                    }),
            .out_data(lut_783_out)
        );

reg   lut_783_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_783_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_783_ff <= lut_783_out;
    end
end

assign out_data[783] = lut_783_ff;




// LUT : 784

wire lut_784_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100010000110111100001000001001110100100000101111010001000000),
            .DEVICE(DEVICE)
        )
    i_lut_784
        (
            .in_data({
                         in_data[434],
                         in_data[520],
                         in_data[557],
                         in_data[76],
                         in_data[506],
                         in_data[403]
                    }),
            .out_data(lut_784_out)
        );

reg   lut_784_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_784_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_784_ff <= lut_784_out;
    end
end

assign out_data[784] = lut_784_ff;




// LUT : 785

wire lut_785_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001001001111010110011110011001000001010111110100011101001101010),
            .DEVICE(DEVICE)
        )
    i_lut_785
        (
            .in_data({
                         in_data[418],
                         in_data[425],
                         in_data[469],
                         in_data[761],
                         in_data[213],
                         in_data[541]
                    }),
            .out_data(lut_785_out)
        );

reg   lut_785_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_785_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_785_ff <= lut_785_out;
    end
end

assign out_data[785] = lut_785_ff;




// LUT : 786

wire lut_786_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011101100100110010111110101100111011111101110001000011010100),
            .DEVICE(DEVICE)
        )
    i_lut_786
        (
            .in_data({
                         in_data[676],
                         in_data[190],
                         in_data[71],
                         in_data[438],
                         in_data[130],
                         in_data[753]
                    }),
            .out_data(lut_786_out)
        );

reg   lut_786_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_786_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_786_ff <= lut_786_out;
    end
end

assign out_data[786] = lut_786_ff;




// LUT : 787

wire lut_787_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100000001110011000011000110011011111100000011000000110100111),
            .DEVICE(DEVICE)
        )
    i_lut_787
        (
            .in_data({
                         in_data[226],
                         in_data[273],
                         in_data[759],
                         in_data[341],
                         in_data[724],
                         in_data[159]
                    }),
            .out_data(lut_787_out)
        );

reg   lut_787_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_787_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_787_ff <= lut_787_out;
    end
end

assign out_data[787] = lut_787_ff;




// LUT : 788

wire lut_788_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010110001110010101000011100000100101111001101001101000111101010),
            .DEVICE(DEVICE)
        )
    i_lut_788
        (
            .in_data({
                         in_data[483],
                         in_data[54],
                         in_data[486],
                         in_data[678],
                         in_data[390],
                         in_data[85]
                    }),
            .out_data(lut_788_out)
        );

reg   lut_788_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_788_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_788_ff <= lut_788_out;
    end
end

assign out_data[788] = lut_788_ff;




// LUT : 789

wire lut_789_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111100010011101111111011111100000110000101111110111011111100),
            .DEVICE(DEVICE)
        )
    i_lut_789
        (
            .in_data({
                         in_data[655],
                         in_data[460],
                         in_data[208],
                         in_data[380],
                         in_data[635],
                         in_data[578]
                    }),
            .out_data(lut_789_out)
        );

reg   lut_789_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_789_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_789_ff <= lut_789_out;
    end
end

assign out_data[789] = lut_789_ff;




// LUT : 790

wire lut_790_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011001011010101001001101000011111010000000001011111000001011),
            .DEVICE(DEVICE)
        )
    i_lut_790
        (
            .in_data({
                         in_data[14],
                         in_data[294],
                         in_data[223],
                         in_data[349],
                         in_data[712],
                         in_data[684]
                    }),
            .out_data(lut_790_out)
        );

reg   lut_790_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_790_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_790_ff <= lut_790_out;
    end
end

assign out_data[790] = lut_790_ff;




// LUT : 791

wire lut_791_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000011001011111011101100110011101011111100110101011111011111),
            .DEVICE(DEVICE)
        )
    i_lut_791
        (
            .in_data({
                         in_data[720],
                         in_data[140],
                         in_data[677],
                         in_data[27],
                         in_data[394],
                         in_data[735]
                    }),
            .out_data(lut_791_out)
        );

reg   lut_791_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_791_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_791_ff <= lut_791_out;
    end
end

assign out_data[791] = lut_791_ff;




// LUT : 792

wire lut_792_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000010000101111011000110000001100110101111111100011111000001),
            .DEVICE(DEVICE)
        )
    i_lut_792
        (
            .in_data({
                         in_data[563],
                         in_data[758],
                         in_data[286],
                         in_data[502],
                         in_data[387],
                         in_data[276]
                    }),
            .out_data(lut_792_out)
        );

reg   lut_792_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_792_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_792_ff <= lut_792_out;
    end
end

assign out_data[792] = lut_792_ff;




// LUT : 793

wire lut_793_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010110011111101110111011101010101110111011101110101111110011010),
            .DEVICE(DEVICE)
        )
    i_lut_793
        (
            .in_data({
                         in_data[499],
                         in_data[135],
                         in_data[611],
                         in_data[428],
                         in_data[302],
                         in_data[778]
                    }),
            .out_data(lut_793_out)
        );

reg   lut_793_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_793_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_793_ff <= lut_793_out;
    end
end

assign out_data[793] = lut_793_ff;




// LUT : 794

wire lut_794_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011010111100010000100101101101001110100000000111101000100010),
            .DEVICE(DEVICE)
        )
    i_lut_794
        (
            .in_data({
                         in_data[24],
                         in_data[311],
                         in_data[112],
                         in_data[391],
                         in_data[429],
                         in_data[455]
                    }),
            .out_data(lut_794_out)
        );

reg   lut_794_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_794_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_794_ff <= lut_794_out;
    end
end

assign out_data[794] = lut_794_ff;




// LUT : 795

wire lut_795_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000010111010000100101100101000011111110010000001000010001000),
            .DEVICE(DEVICE)
        )
    i_lut_795
        (
            .in_data({
                         in_data[30],
                         in_data[439],
                         in_data[84],
                         in_data[480],
                         in_data[315],
                         in_data[13]
                    }),
            .out_data(lut_795_out)
        );

reg   lut_795_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_795_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_795_ff <= lut_795_out;
    end
end

assign out_data[795] = lut_795_ff;




// LUT : 796

wire lut_796_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100111010011011111011110111101010011101011110101111001010101),
            .DEVICE(DEVICE)
        )
    i_lut_796
        (
            .in_data({
                         in_data[309],
                         in_data[612],
                         in_data[229],
                         in_data[703],
                         in_data[437],
                         in_data[123]
                    }),
            .out_data(lut_796_out)
        );

reg   lut_796_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_796_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_796_ff <= lut_796_out;
    end
end

assign out_data[796] = lut_796_ff;




// LUT : 797

wire lut_797_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101101001000001101101100111000001011010010101101010000001010),
            .DEVICE(DEVICE)
        )
    i_lut_797
        (
            .in_data({
                         in_data[269],
                         in_data[161],
                         in_data[743],
                         in_data[136],
                         in_data[535],
                         in_data[651]
                    }),
            .out_data(lut_797_out)
        );

reg   lut_797_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_797_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_797_ff <= lut_797_out;
    end
end

assign out_data[797] = lut_797_ff;




// LUT : 798

wire lut_798_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101111111010110011001001100011000111011000111101000011011110),
            .DEVICE(DEVICE)
        )
    i_lut_798
        (
            .in_data({
                         in_data[266],
                         in_data[306],
                         in_data[262],
                         in_data[322],
                         in_data[285],
                         in_data[316]
                    }),
            .out_data(lut_798_out)
        );

reg   lut_798_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_798_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_798_ff <= lut_798_out;
    end
end

assign out_data[798] = lut_798_ff;




// LUT : 799

wire lut_799_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100001100111001000101110111010100101011100101110110110101011100),
            .DEVICE(DEVICE)
        )
    i_lut_799
        (
            .in_data({
                         in_data[171],
                         in_data[228],
                         in_data[622],
                         in_data[128],
                         in_data[141],
                         in_data[443]
                    }),
            .out_data(lut_799_out)
        );

reg   lut_799_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_799_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_799_ff <= lut_799_out;
    end
end

assign out_data[799] = lut_799_ff;




// LUT : 800

wire lut_800_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100110111111100100101101100110100111000101011101001110111101),
            .DEVICE(DEVICE)
        )
    i_lut_800
        (
            .in_data({
                         in_data[82],
                         in_data[156],
                         in_data[771],
                         in_data[290],
                         in_data[3],
                         in_data[644]
                    }),
            .out_data(lut_800_out)
        );

reg   lut_800_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_800_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_800_ff <= lut_800_out;
    end
end

assign out_data[800] = lut_800_ff;




// LUT : 801

wire lut_801_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111100010110101111101100111011011101101011110010111111010101010),
            .DEVICE(DEVICE)
        )
    i_lut_801
        (
            .in_data({
                         in_data[625],
                         in_data[531],
                         in_data[683],
                         in_data[544],
                         in_data[230],
                         in_data[92]
                    }),
            .out_data(lut_801_out)
        );

reg   lut_801_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_801_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_801_ff <= lut_801_out;
    end
end

assign out_data[801] = lut_801_ff;




// LUT : 802

wire lut_802_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101010111001111000000000000010100000001000000000010010100100),
            .DEVICE(DEVICE)
        )
    i_lut_802
        (
            .in_data({
                         in_data[479],
                         in_data[324],
                         in_data[685],
                         in_data[166],
                         in_data[410],
                         in_data[621]
                    }),
            .out_data(lut_802_out)
        );

reg   lut_802_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_802_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_802_ff <= lut_802_out;
    end
end

assign out_data[802] = lut_802_ff;




// LUT : 803

wire lut_803_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111010111110101110001111000001101010010011000000100010001010),
            .DEVICE(DEVICE)
        )
    i_lut_803
        (
            .in_data({
                         in_data[649],
                         in_data[670],
                         in_data[601],
                         in_data[250],
                         in_data[664],
                         in_data[323]
                    }),
            .out_data(lut_803_out)
        );

reg   lut_803_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_803_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_803_ff <= lut_803_out;
    end
end

assign out_data[803] = lut_803_ff;




// LUT : 804

wire lut_804_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001110000110000010011000001000001001111111100000000011111010001),
            .DEVICE(DEVICE)
        )
    i_lut_804
        (
            .in_data({
                         in_data[371],
                         in_data[291],
                         in_data[476],
                         in_data[86],
                         in_data[546],
                         in_data[426]
                    }),
            .out_data(lut_804_out)
        );

reg   lut_804_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_804_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_804_ff <= lut_804_out;
    end
end

assign out_data[804] = lut_804_ff;




// LUT : 805

wire lut_805_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011001001100010010010100101011011101101000101101111000001010),
            .DEVICE(DEVICE)
        )
    i_lut_805
        (
            .in_data({
                         in_data[490],
                         in_data[67],
                         in_data[16],
                         in_data[393],
                         in_data[717],
                         in_data[628]
                    }),
            .out_data(lut_805_out)
        );

reg   lut_805_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_805_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_805_ff <= lut_805_out;
    end
end

assign out_data[805] = lut_805_ff;




// LUT : 806

wire lut_806_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001100001111010001011101001110010101010111011010000011101000010),
            .DEVICE(DEVICE)
        )
    i_lut_806
        (
            .in_data({
                         in_data[210],
                         in_data[53],
                         in_data[591],
                         in_data[8],
                         in_data[671],
                         in_data[150]
                    }),
            .out_data(lut_806_out)
        );

reg   lut_806_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_806_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_806_ff <= lut_806_out;
    end
end

assign out_data[806] = lut_806_ff;




// LUT : 807

wire lut_807_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111111111111001010101010101010111111111111110000100000001000),
            .DEVICE(DEVICE)
        )
    i_lut_807
        (
            .in_data({
                         in_data[217],
                         in_data[408],
                         in_data[414],
                         in_data[398],
                         in_data[244],
                         in_data[451]
                    }),
            .out_data(lut_807_out)
        );

reg   lut_807_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_807_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_807_ff <= lut_807_out;
    end
end

assign out_data[807] = lut_807_ff;




// LUT : 808

wire lut_808_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010110000100010000010000000101011111100010010100000100000000),
            .DEVICE(DEVICE)
        )
    i_lut_808
        (
            .in_data({
                         in_data[180],
                         in_data[293],
                         in_data[234],
                         in_data[584],
                         in_data[399],
                         in_data[609]
                    }),
            .out_data(lut_808_out)
        );

reg   lut_808_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_808_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_808_ff <= lut_808_out;
    end
end

assign out_data[808] = lut_808_ff;




// LUT : 809

wire lut_809_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000001001000011001100001000000001001101110010000100110001001),
            .DEVICE(DEVICE)
        )
    i_lut_809
        (
            .in_data({
                         in_data[705],
                         in_data[627],
                         in_data[608],
                         in_data[218],
                         in_data[507],
                         in_data[219]
                    }),
            .out_data(lut_809_out)
        );

reg   lut_809_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_809_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_809_ff <= lut_809_out;
    end
end

assign out_data[809] = lut_809_ff;




// LUT : 810

wire lut_810_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101011001111110000101100110100101101100111000101001000011001),
            .DEVICE(DEVICE)
        )
    i_lut_810
        (
            .in_data({
                         in_data[132],
                         in_data[533],
                         in_data[253],
                         in_data[109],
                         in_data[767],
                         in_data[81]
                    }),
            .out_data(lut_810_out)
        );

reg   lut_810_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_810_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_810_ff <= lut_810_out;
    end
end

assign out_data[810] = lut_810_ff;




// LUT : 811

wire lut_811_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010010100001100110001011100101110101010001100000101011111101110),
            .DEVICE(DEVICE)
        )
    i_lut_811
        (
            .in_data({
                         in_data[255],
                         in_data[107],
                         in_data[475],
                         in_data[158],
                         in_data[98],
                         in_data[126]
                    }),
            .out_data(lut_811_out)
        );

reg   lut_811_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_811_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_811_ff <= lut_811_out;
    end
end

assign out_data[811] = lut_811_ff;




// LUT : 812

wire lut_812_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001000010000001010101111000010100010000100001111110111010100),
            .DEVICE(DEVICE)
        )
    i_lut_812
        (
            .in_data({
                         in_data[545],
                         in_data[543],
                         in_data[657],
                         in_data[245],
                         in_data[182],
                         in_data[64]
                    }),
            .out_data(lut_812_out)
        );

reg   lut_812_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_812_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_812_ff <= lut_812_out;
    end
end

assign out_data[812] = lut_812_ff;




// LUT : 813

wire lut_813_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001001001001010011110001011110010110100001101101111101101101010),
            .DEVICE(DEVICE)
        )
    i_lut_813
        (
            .in_data({
                         in_data[650],
                         in_data[254],
                         in_data[247],
                         in_data[556],
                         in_data[252],
                         in_data[175]
                    }),
            .out_data(lut_813_out)
        );

reg   lut_813_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_813_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_813_ff <= lut_813_out;
    end
end

assign out_data[813] = lut_813_ff;




// LUT : 814

wire lut_814_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011111111111000101000111010110001100110101111101110110101100),
            .DEVICE(DEVICE)
        )
    i_lut_814
        (
            .in_data({
                         in_data[737],
                         in_data[199],
                         in_data[91],
                         in_data[456],
                         in_data[257],
                         in_data[477]
                    }),
            .out_data(lut_814_out)
        );

reg   lut_814_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_814_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_814_ff <= lut_814_out;
    end
end

assign out_data[814] = lut_814_ff;




// LUT : 815

wire lut_815_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111011101001110000001100101010110010110111000000010001101111),
            .DEVICE(DEVICE)
        )
    i_lut_815
        (
            .in_data({
                         in_data[573],
                         in_data[726],
                         in_data[145],
                         in_data[504],
                         in_data[280],
                         in_data[261]
                    }),
            .out_data(lut_815_out)
        );

reg   lut_815_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_815_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_815_ff <= lut_815_out;
    end
end

assign out_data[815] = lut_815_ff;




// LUT : 816

wire lut_816_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010001100000011100000001110101010000101110001000100011110101),
            .DEVICE(DEVICE)
        )
    i_lut_816
        (
            .in_data({
                         in_data[212],
                         in_data[68],
                         in_data[523],
                         in_data[11],
                         in_data[304],
                         in_data[647]
                    }),
            .out_data(lut_816_out)
        );

reg   lut_816_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_816_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_816_ff <= lut_816_out;
    end
end

assign out_data[816] = lut_816_ff;




// LUT : 817

wire lut_817_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110011000100110010101011000001111101000001110000110010001111110),
            .DEVICE(DEVICE)
        )
    i_lut_817
        (
            .in_data({
                         in_data[746],
                         in_data[623],
                         in_data[231],
                         in_data[447],
                         in_data[139],
                         in_data[605]
                    }),
            .out_data(lut_817_out)
        );

reg   lut_817_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_817_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_817_ff <= lut_817_out;
    end
end

assign out_data[817] = lut_817_ff;




// LUT : 818

wire lut_818_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001010100011011000110110000001001010101111000010100010000101),
            .DEVICE(DEVICE)
        )
    i_lut_818
        (
            .in_data({
                         in_data[15],
                         in_data[144],
                         in_data[339],
                         in_data[74],
                         in_data[146],
                         in_data[590]
                    }),
            .out_data(lut_818_out)
        );

reg   lut_818_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_818_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_818_ff <= lut_818_out;
    end
end

assign out_data[818] = lut_818_ff;




// LUT : 819

wire lut_819_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100010111110101100101011010011011101110101010100111101100000),
            .DEVICE(DEVICE)
        )
    i_lut_819
        (
            .in_data({
                         in_data[752],
                         in_data[292],
                         in_data[312],
                         in_data[423],
                         in_data[400],
                         in_data[404]
                    }),
            .out_data(lut_819_out)
        );

reg   lut_819_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_819_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_819_ff <= lut_819_out;
    end
end

assign out_data[819] = lut_819_ff;




// LUT : 820

wire lut_820_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001000001100111010100010110000001100000110000100010000011001),
            .DEVICE(DEVICE)
        )
    i_lut_820
        (
            .in_data({
                         in_data[589],
                         in_data[610],
                         in_data[133],
                         in_data[656],
                         in_data[747],
                         in_data[177]
                    }),
            .out_data(lut_820_out)
        );

reg   lut_820_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_820_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_820_ff <= lut_820_out;
    end
end

assign out_data[820] = lut_820_ff;




// LUT : 821

wire lut_821_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111101010010110111001010000011110111101000110001000000000001),
            .DEVICE(DEVICE)
        )
    i_lut_821
        (
            .in_data({
                         in_data[221],
                         in_data[666],
                         in_data[618],
                         in_data[689],
                         in_data[631],
                         in_data[94]
                    }),
            .out_data(lut_821_out)
        );

reg   lut_821_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_821_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_821_ff <= lut_821_out;
    end
end

assign out_data[821] = lut_821_ff;




// LUT : 822

wire lut_822_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110110010110110101100001101011100010101111001011100111100010011),
            .DEVICE(DEVICE)
        )
    i_lut_822
        (
            .in_data({
                         in_data[51],
                         in_data[662],
                         in_data[348],
                         in_data[364],
                         in_data[205],
                         in_data[653]
                    }),
            .out_data(lut_822_out)
        );

reg   lut_822_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_822_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_822_ff <= lut_822_out;
    end
end

assign out_data[822] = lut_822_ff;




// LUT : 823

wire lut_823_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010010100011001111101011010001101111011100010111101011001100),
            .DEVICE(DEVICE)
        )
    i_lut_823
        (
            .in_data({
                         in_data[588],
                         in_data[736],
                         in_data[757],
                         in_data[232],
                         in_data[714],
                         in_data[532]
                    }),
            .out_data(lut_823_out)
        );

reg   lut_823_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_823_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_823_ff <= lut_823_out;
    end
end

assign out_data[823] = lut_823_ff;




// LUT : 824

wire lut_824_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110011001000000111100000111101001000000111011111010011101101111),
            .DEVICE(DEVICE)
        )
    i_lut_824
        (
            .in_data({
                         in_data[774],
                         in_data[687],
                         in_data[289],
                         in_data[164],
                         in_data[478],
                         in_data[89]
                    }),
            .out_data(lut_824_out)
        );

reg   lut_824_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_824_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_824_ff <= lut_824_out;
    end
end

assign out_data[824] = lut_824_ff;




// LUT : 825

wire lut_825_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100010011001101101000111111111001111011000110000110110111011),
            .DEVICE(DEVICE)
        )
    i_lut_825
        (
            .in_data({
                         in_data[87],
                         in_data[56],
                         in_data[643],
                         in_data[780],
                         in_data[376],
                         in_data[615]
                    }),
            .out_data(lut_825_out)
        );

reg   lut_825_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_825_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_825_ff <= lut_825_out;
    end
end

assign out_data[825] = lut_825_ff;




// LUT : 826

wire lut_826_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111111001100111100010101010111111111010101011100000010011100),
            .DEVICE(DEVICE)
        )
    i_lut_826
        (
            .in_data({
                         in_data[763],
                         in_data[472],
                         in_data[467],
                         in_data[327],
                         in_data[19],
                         in_data[660]
                    }),
            .out_data(lut_826_out)
        );

reg   lut_826_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_826_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_826_ff <= lut_826_out;
    end
end

assign out_data[826] = lut_826_ff;




// LUT : 827

wire lut_827_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001001110011101010111110111100110101111101011111100011111100111),
            .DEVICE(DEVICE)
        )
    i_lut_827
        (
            .in_data({
                         in_data[783],
                         in_data[512],
                         in_data[272],
                         in_data[235],
                         in_data[554],
                         in_data[101]
                    }),
            .out_data(lut_827_out)
        );

reg   lut_827_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_827_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_827_ff <= lut_827_out;
    end
end

assign out_data[827] = lut_827_ff;




// LUT : 828

wire lut_828_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001001000010110000011000110101001000010111001011110010101100),
            .DEVICE(DEVICE)
        )
    i_lut_828
        (
            .in_data({
                         in_data[365],
                         in_data[153],
                         in_data[526],
                         in_data[673],
                         in_data[482],
                         in_data[242]
                    }),
            .out_data(lut_828_out)
        );

reg   lut_828_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_828_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_828_ff <= lut_828_out;
    end
end

assign out_data[828] = lut_828_ff;




// LUT : 829

wire lut_829_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110011110111001001010000011111001111100011010001111000011010101),
            .DEVICE(DEVICE)
        )
    i_lut_829
        (
            .in_data({
                         in_data[688],
                         in_data[674],
                         in_data[494],
                         in_data[196],
                         in_data[412],
                         in_data[121]
                    }),
            .out_data(lut_829_out)
        );

reg   lut_829_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_829_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_829_ff <= lut_829_out;
    end
end

assign out_data[829] = lut_829_ff;




// LUT : 830

wire lut_830_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000100000101010111000101111111011110111111110011100001001110),
            .DEVICE(DEVICE)
        )
    i_lut_830
        (
            .in_data({
                         in_data[637],
                         in_data[39],
                         in_data[755],
                         in_data[381],
                         in_data[149],
                         in_data[385]
                    }),
            .out_data(lut_830_out)
        );

reg   lut_830_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_830_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_830_ff <= lut_830_out;
    end
end

assign out_data[830] = lut_830_ff;




// LUT : 831

wire lut_831_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001001100010011001101010110110001000110001011110101000001001),
            .DEVICE(DEVICE)
        )
    i_lut_831
        (
            .in_data({
                         in_data[360],
                         in_data[754],
                         in_data[114],
                         in_data[186],
                         in_data[421],
                         in_data[730]
                    }),
            .out_data(lut_831_out)
        );

reg   lut_831_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_831_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_831_ff <= lut_831_out;
    end
end

assign out_data[831] = lut_831_ff;




// LUT : 832

wire lut_832_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100010101011011101000100010000011100110111001110100010100000),
            .DEVICE(DEVICE)
        )
    i_lut_832
        (
            .in_data({
                         in_data[595],
                         in_data[699],
                         in_data[681],
                         in_data[201],
                         in_data[407],
                         in_data[484]
                    }),
            .out_data(lut_832_out)
        );

reg   lut_832_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_832_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_832_ff <= lut_832_out;
    end
end

assign out_data[832] = lut_832_ff;




// LUT : 833

wire lut_833_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101101110101100000100000001100011000000000000000000010100001101),
            .DEVICE(DEVICE)
        )
    i_lut_833
        (
            .in_data({
                         in_data[78],
                         in_data[120],
                         in_data[440],
                         in_data[632],
                         in_data[246],
                         in_data[540]
                    }),
            .out_data(lut_833_out)
        );

reg   lut_833_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_833_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_833_ff <= lut_833_out;
    end
end

assign out_data[833] = lut_833_ff;




// LUT : 834

wire lut_834_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001000111100110100000000000101101101100000001010000000100001),
            .DEVICE(DEVICE)
        )
    i_lut_834
        (
            .in_data({
                         in_data[417],
                         in_data[503],
                         in_data[734],
                         in_data[581],
                         in_data[716],
                         in_data[331]
                    }),
            .out_data(lut_834_out)
        );

reg   lut_834_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_834_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_834_ff <= lut_834_out;
    end
end

assign out_data[834] = lut_834_ff;




// LUT : 835

wire lut_835_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110000011110000000010101001110010100010101000000110110100001),
            .DEVICE(DEVICE)
        )
    i_lut_835
        (
            .in_data({
                         in_data[137],
                         in_data[36],
                         in_data[654],
                         in_data[382],
                         in_data[413],
                         in_data[619]
                    }),
            .out_data(lut_835_out)
        );

reg   lut_835_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_835_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_835_ff <= lut_835_out;
    end
end

assign out_data[835] = lut_835_ff;




// LUT : 836

wire lut_836_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100010111101001001010001011111010010100100001100101010010001),
            .DEVICE(DEVICE)
        )
    i_lut_836
        (
            .in_data({
                         in_data[191],
                         in_data[713],
                         in_data[667],
                         in_data[192],
                         in_data[359],
                         in_data[63]
                    }),
            .out_data(lut_836_out)
        );

reg   lut_836_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_836_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_836_ff <= lut_836_out;
    end
end

assign out_data[836] = lut_836_ff;




// LUT : 837

wire lut_837_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100001010011010110101011111010011010111010100011111111101110011),
            .DEVICE(DEVICE)
        )
    i_lut_837
        (
            .in_data({
                         in_data[181],
                         in_data[765],
                         in_data[305],
                         in_data[372],
                         in_data[492],
                         in_data[227]
                    }),
            .out_data(lut_837_out)
        );

reg   lut_837_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_837_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_837_ff <= lut_837_out;
    end
end

assign out_data[837] = lut_837_ff;




// LUT : 838

wire lut_838_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100100100101000011101111111111111010101011001111100011111101),
            .DEVICE(DEVICE)
        )
    i_lut_838
        (
            .in_data({
                         in_data[9],
                         in_data[441],
                         in_data[263],
                         in_data[310],
                         in_data[202],
                         in_data[715]
                    }),
            .out_data(lut_838_out)
        );

reg   lut_838_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_838_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_838_ff <= lut_838_out;
    end
end

assign out_data[838] = lut_838_ff;




// LUT : 839

wire lut_839_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111101001001100100011001001110000101100010101001011111001000011),
            .DEVICE(DEVICE)
        )
    i_lut_839
        (
            .in_data({
                         in_data[313],
                         in_data[62],
                         in_data[663],
                         in_data[629],
                         in_data[45],
                         in_data[301]
                    }),
            .out_data(lut_839_out)
        );

reg   lut_839_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_839_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_839_ff <= lut_839_out;
    end
end

assign out_data[839] = lut_839_ff;




// LUT : 840

wire lut_840_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110011000100000110111101011100101100010101100011101110000111101),
            .DEVICE(DEVICE)
        )
    i_lut_840
        (
            .in_data({
                         in_data[179],
                         in_data[491],
                         in_data[106],
                         in_data[593],
                         in_data[115],
                         in_data[277]
                    }),
            .out_data(lut_840_out)
        );

reg   lut_840_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_840_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_840_ff <= lut_840_out;
    end
end

assign out_data[840] = lut_840_ff;




// LUT : 841

wire lut_841_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010111110110100001000000110100011101100011000000111101011001),
            .DEVICE(DEVICE)
        )
    i_lut_841
        (
            .in_data({
                         in_data[185],
                         in_data[4],
                         in_data[251],
                         in_data[134],
                         in_data[275],
                         in_data[411]
                    }),
            .out_data(lut_841_out)
        );

reg   lut_841_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_841_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_841_ff <= lut_841_out;
    end
end

assign out_data[841] = lut_841_ff;




// LUT : 842

wire lut_842_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111100100010101101011110111011110100111011101010000110111010100),
            .DEVICE(DEVICE)
        )
    i_lut_842
        (
            .in_data({
                         in_data[522],
                         in_data[594],
                         in_data[587],
                         in_data[93],
                         in_data[165],
                         in_data[7]
                    }),
            .out_data(lut_842_out)
        );

reg   lut_842_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_842_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_842_ff <= lut_842_out;
    end
end

assign out_data[842] = lut_842_ff;




// LUT : 843

wire lut_843_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001001101010100101001111100111010110010111011000011011111110),
            .DEVICE(DEVICE)
        )
    i_lut_843
        (
            .in_data({
                         in_data[358],
                         in_data[583],
                         in_data[749],
                         in_data[596],
                         in_data[97],
                         in_data[18]
                    }),
            .out_data(lut_843_out)
        );

reg   lut_843_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_843_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_843_ff <= lut_843_out;
    end
end

assign out_data[843] = lut_843_ff;




// LUT : 844

wire lut_844_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000010110110000011111111111110111111010001001011111100101000),
            .DEVICE(DEVICE)
        )
    i_lut_844
        (
            .in_data({
                         in_data[680],
                         in_data[129],
                         in_data[693],
                         in_data[462],
                         in_data[189],
                         in_data[727]
                    }),
            .out_data(lut_844_out)
        );

reg   lut_844_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_844_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_844_ff <= lut_844_out;
    end
end

assign out_data[844] = lut_844_ff;




// LUT : 845

wire lut_845_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101111101011110010111010111010111111111000101110000011001100),
            .DEVICE(DEVICE)
        )
    i_lut_845
        (
            .in_data({
                         in_data[26],
                         in_data[334],
                         in_data[25],
                         in_data[464],
                         in_data[745],
                         in_data[342]
                    }),
            .out_data(lut_845_out)
        );

reg   lut_845_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_845_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_845_ff <= lut_845_out;
    end
end

assign out_data[845] = lut_845_ff;




// LUT : 846

wire lut_846_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010101100101011000000011111110000010101110101100101111000001),
            .DEVICE(DEVICE)
        )
    i_lut_846
        (
            .in_data({
                         in_data[766],
                         in_data[518],
                         in_data[238],
                         in_data[57],
                         in_data[640],
                         in_data[560]
                    }),
            .out_data(lut_846_out)
        );

reg   lut_846_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_846_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_846_ff <= lut_846_out;
    end
end

assign out_data[846] = lut_846_ff;




// LUT : 847

wire lut_847_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101011010101001101100001111010000101111110111111111111110110),
            .DEVICE(DEVICE)
        )
    i_lut_847
        (
            .in_data({
                         in_data[652],
                         in_data[524],
                         in_data[102],
                         in_data[268],
                         in_data[592],
                         in_data[113]
                    }),
            .out_data(lut_847_out)
        );

reg   lut_847_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_847_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_847_ff <= lut_847_out;
    end
end

assign out_data[847] = lut_847_ff;




// LUT : 848

wire lut_848_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000100101001111010001110100000110111111001101001001101010011),
            .DEVICE(DEVICE)
        )
    i_lut_848
        (
            .in_data({
                         in_data[222],
                         in_data[682],
                         in_data[206],
                         in_data[728],
                         in_data[772],
                         in_data[579]
                    }),
            .out_data(lut_848_out)
        );

reg   lut_848_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_848_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_848_ff <= lut_848_out;
    end
end

assign out_data[848] = lut_848_ff;




// LUT : 849

wire lut_849_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001101101110101011001000110001001000000000100100000000000001),
            .DEVICE(DEVICE)
        )
    i_lut_849
        (
            .in_data({
                         in_data[698],
                         in_data[549],
                         in_data[77],
                         in_data[386],
                         in_data[770],
                         in_data[602]
                    }),
            .out_data(lut_849_out)
        );

reg   lut_849_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_849_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_849_ff <= lut_849_out;
    end
end

assign out_data[849] = lut_849_ff;




// LUT : 850

wire lut_850_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000110110110100111001110111100001011010101101011010111010110),
            .DEVICE(DEVICE)
        )
    i_lut_850
        (
            .in_data({
                         in_data[154],
                         in_data[168],
                         in_data[762],
                         in_data[642],
                         in_data[328],
                         in_data[598]
                    }),
            .out_data(lut_850_out)
        );

reg   lut_850_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_850_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_850_ff <= lut_850_out;
    end
end

assign out_data[850] = lut_850_ff;




// LUT : 851

wire lut_851_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111011001000101011000111110111000100101010111101011100110011),
            .DEVICE(DEVICE)
        )
    i_lut_851
        (
            .in_data({
                         in_data[340],
                         in_data[599],
                         in_data[49],
                         in_data[686],
                         in_data[442],
                         in_data[646]
                    }),
            .out_data(lut_851_out)
        );

reg   lut_851_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_851_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_851_ff <= lut_851_out;
    end
end

assign out_data[851] = lut_851_ff;




// LUT : 852

wire lut_852_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110111001100000011101111111100011111111010110100000111100011000),
            .DEVICE(DEVICE)
        )
    i_lut_852
        (
            .in_data({
                         in_data[66],
                         in_data[216],
                         in_data[537],
                         in_data[264],
                         in_data[466],
                         in_data[634]
                    }),
            .out_data(lut_852_out)
        );

reg   lut_852_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_852_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_852_ff <= lut_852_out;
    end
end

assign out_data[852] = lut_852_ff;




// LUT : 853

wire lut_853_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110110101001100010010110101011111101101111111101111111111010),
            .DEVICE(DEVICE)
        )
    i_lut_853
        (
            .in_data({
                         in_data[237],
                         in_data[748],
                         in_data[42],
                         in_data[1],
                         in_data[433],
                         in_data[487]
                    }),
            .out_data(lut_853_out)
        );

reg   lut_853_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_853_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_853_ff <= lut_853_out;
    end
end

assign out_data[853] = lut_853_ff;




// LUT : 854

wire lut_854_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001100101000001110010111101110101100110010000100100100101110),
            .DEVICE(DEVICE)
        )
    i_lut_854
        (
            .in_data({
                         in_data[178],
                         in_data[155],
                         in_data[40],
                         in_data[641],
                         in_data[103],
                         in_data[694]
                    }),
            .out_data(lut_854_out)
        );

reg   lut_854_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_854_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_854_ff <= lut_854_out;
    end
end

assign out_data[854] = lut_854_ff;




// LUT : 855

wire lut_855_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010110001011100111111111100010110011101110110010110011111111),
            .DEVICE(DEVICE)
        )
    i_lut_855
        (
            .in_data({
                         in_data[281],
                         in_data[706],
                         in_data[569],
                         in_data[431],
                         in_data[124],
                         in_data[567]
                    }),
            .out_data(lut_855_out)
        );

reg   lut_855_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_855_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_855_ff <= lut_855_out;
    end
end

assign out_data[855] = lut_855_ff;




// LUT : 856

wire lut_856_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111100100100110100110101011110010111100000000100101000010000),
            .DEVICE(DEVICE)
        )
    i_lut_856
        (
            .in_data({
                         in_data[461],
                         in_data[675],
                         in_data[127],
                         in_data[719],
                         in_data[709],
                         in_data[353]
                    }),
            .out_data(lut_856_out)
        );

reg   lut_856_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_856_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_856_ff <= lut_856_out;
    end
end

assign out_data[856] = lut_856_ff;




// LUT : 857

wire lut_857_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111001001111110110000011000100100110000000010110000011111101),
            .DEVICE(DEVICE)
        )
    i_lut_857
        (
            .in_data({
                         in_data[459],
                         in_data[711],
                         in_data[256],
                         in_data[616],
                         in_data[17],
                         in_data[197]
                    }),
            .out_data(lut_857_out)
        );

reg   lut_857_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_857_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_857_ff <= lut_857_out;
    end
end

assign out_data[857] = lut_857_ff;




// LUT : 858

wire lut_858_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010110100101111111111011111010001100111111111010001100100011),
            .DEVICE(DEVICE)
        )
    i_lut_858
        (
            .in_data({
                         in_data[528],
                         in_data[722],
                         in_data[513],
                         in_data[183],
                         in_data[233],
                         in_data[240]
                    }),
            .out_data(lut_858_out)
        );

reg   lut_858_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_858_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_858_ff <= lut_858_out;
    end
end

assign out_data[858] = lut_858_ff;




// LUT : 859

wire lut_859_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001001010001110011111000101001110111001101011101011101101100110),
            .DEVICE(DEVICE)
        )
    i_lut_859
        (
            .in_data({
                         in_data[279],
                         in_data[314],
                         in_data[95],
                         in_data[539],
                         in_data[138],
                         in_data[152]
                    }),
            .out_data(lut_859_out)
        );

reg   lut_859_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_859_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_859_ff <= lut_859_out;
    end
end

assign out_data[859] = lut_859_ff;




// LUT : 860

wire lut_860_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110100110010010100011001111111100110000111100111111111110101),
            .DEVICE(DEVICE)
        )
    i_lut_860
        (
            .in_data({
                         in_data[718],
                         in_data[782],
                         in_data[561],
                         in_data[739],
                         in_data[457],
                         in_data[525]
                    }),
            .out_data(lut_860_out)
        );

reg   lut_860_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_860_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_860_ff <= lut_860_out;
    end
end

assign out_data[860] = lut_860_ff;




// LUT : 861

wire lut_861_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111110001111010111110110111010100000111011000011001111101011),
            .DEVICE(DEVICE)
        )
    i_lut_861
        (
            .in_data({
                         in_data[721],
                         in_data[329],
                         in_data[401],
                         in_data[147],
                         in_data[355],
                         in_data[468]
                    }),
            .out_data(lut_861_out)
        );

reg   lut_861_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_861_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_861_ff <= lut_861_out;
    end
end

assign out_data[861] = lut_861_ff;




// LUT : 862

wire lut_862_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100101111110110000101000001101111111000000001011001110110010),
            .DEVICE(DEVICE)
        )
    i_lut_862
        (
            .in_data({
                         in_data[308],
                         in_data[529],
                         in_data[288],
                         in_data[550],
                         in_data[295],
                         in_data[430]
                    }),
            .out_data(lut_862_out)
        );

reg   lut_862_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_862_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_862_ff <= lut_862_out;
    end
end

assign out_data[862] = lut_862_ff;




// LUT : 863

wire lut_863_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100100001000001011010111111011000100010101000011001100110000),
            .DEVICE(DEVICE)
        )
    i_lut_863
        (
            .in_data({
                         in_data[282],
                         in_data[105],
                         in_data[248],
                         in_data[363],
                         in_data[37],
                         in_data[542]
                    }),
            .out_data(lut_863_out)
        );

reg   lut_863_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_863_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_863_ff <= lut_863_out;
    end
end

assign out_data[863] = lut_863_ff;




// LUT : 864

wire lut_864_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010001001000100010100100110100010110000011000110110100000001),
            .DEVICE(DEVICE)
        )
    i_lut_864
        (
            .in_data({
                         in_data[445],
                         in_data[69],
                         in_data[530],
                         in_data[501],
                         in_data[725],
                         in_data[572]
                    }),
            .out_data(lut_864_out)
        );

reg   lut_864_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_864_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_864_ff <= lut_864_out;
    end
end

assign out_data[864] = lut_864_ff;




// LUT : 865

wire lut_865_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101101101110110010010111001101010110111011101111101101111111),
            .DEVICE(DEVICE)
        )
    i_lut_865
        (
            .in_data({
                         in_data[565],
                         in_data[35],
                         in_data[750],
                         in_data[744],
                         in_data[303],
                         in_data[775]
                    }),
            .out_data(lut_865_out)
        );

reg   lut_865_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_865_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_865_ff <= lut_865_out;
    end
end

assign out_data[865] = lut_865_ff;




// LUT : 866

wire lut_866_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011100000001000111110001000010100111001111111111011101110001),
            .DEVICE(DEVICE)
        )
    i_lut_866
        (
            .in_data({
                         in_data[214],
                         in_data[639],
                         in_data[270],
                         in_data[695],
                         in_data[638],
                         in_data[626]
                    }),
            .out_data(lut_866_out)
        );

reg   lut_866_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_866_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_866_ff <= lut_866_out;
    end
end

assign out_data[866] = lut_866_ff;




// LUT : 867

wire lut_867_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011100001001101011110001011111000010000000001011110100000001),
            .DEVICE(DEVICE)
        )
    i_lut_867
        (
            .in_data({
                         in_data[769],
                         in_data[160],
                         in_data[760],
                         in_data[521],
                         in_data[204],
                         in_data[187]
                    }),
            .out_data(lut_867_out)
        );

reg   lut_867_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_867_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_867_ff <= lut_867_out;
    end
end

assign out_data[867] = lut_867_ff;




// LUT : 868

wire lut_868_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111101000111001010011010000110000010011001101011111111101011101),
            .DEVICE(DEVICE)
        )
    i_lut_868
        (
            .in_data({
                         in_data[243],
                         in_data[29],
                         in_data[357],
                         in_data[298],
                         in_data[516],
                         in_data[347]
                    }),
            .out_data(lut_868_out)
        );

reg   lut_868_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_868_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_868_ff <= lut_868_out;
    end
end

assign out_data[868] = lut_868_ff;




// LUT : 869

wire lut_869_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101001011010111100111100111111000001111011111000001101001011110),
            .DEVICE(DEVICE)
        )
    i_lut_869
        (
            .in_data({
                         in_data[297],
                         in_data[283],
                         in_data[117],
                         in_data[259],
                         in_data[741],
                         in_data[23]
                    }),
            .out_data(lut_869_out)
        );

reg   lut_869_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_869_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_869_ff <= lut_869_out;
    end
end

assign out_data[869] = lut_869_ff;




// LUT : 870

wire lut_870_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000011111101110010000101010001101000111110111001110000000001),
            .DEVICE(DEVICE)
        )
    i_lut_870
        (
            .in_data({
                         in_data[493],
                         in_data[296],
                         in_data[648],
                         in_data[96],
                         in_data[148],
                         in_data[354]
                    }),
            .out_data(lut_870_out)
        );

reg   lut_870_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_870_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_870_ff <= lut_870_out;
    end
end

assign out_data[870] = lut_870_ff;




// LUT : 871

wire lut_871_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000000000000010100010000000010011110101100011101110010100101),
            .DEVICE(DEVICE)
        )
    i_lut_871
        (
            .in_data({
                         in_data[510],
                         in_data[267],
                         in_data[474],
                         in_data[20],
                         in_data[564],
                         in_data[452]
                    }),
            .out_data(lut_871_out)
        );

reg   lut_871_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_871_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_871_ff <= lut_871_out;
    end
end

assign out_data[871] = lut_871_ff;




// LUT : 872

wire lut_872_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111101110011101101111110010110111101011011110101011101101010),
            .DEVICE(DEVICE)
        )
    i_lut_872
        (
            .in_data({
                         in_data[351],
                         in_data[325],
                         in_data[90],
                         in_data[370],
                         in_data[28],
                         in_data[751]
                    }),
            .out_data(lut_872_out)
        );

reg   lut_872_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_872_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_872_ff <= lut_872_out;
    end
end

assign out_data[872] = lut_872_ff;




// LUT : 873

wire lut_873_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010100000000000011010000100101000000110110001100000011111001),
            .DEVICE(DEVICE)
        )
    i_lut_873
        (
            .in_data({
                         in_data[388],
                         in_data[435],
                         in_data[125],
                         in_data[630],
                         in_data[317],
                         in_data[661]
                    }),
            .out_data(lut_873_out)
        );

reg   lut_873_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_873_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_873_ff <= lut_873_out;
    end
end

assign out_data[873] = lut_873_ff;




// LUT : 874

wire lut_874_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101000001010111100111110010000000011100010001110111111101001),
            .DEVICE(DEVICE)
        )
    i_lut_874
        (
            .in_data({
                         in_data[489],
                         in_data[207],
                         in_data[321],
                         in_data[568],
                         in_data[415],
                         in_data[781]
                    }),
            .out_data(lut_874_out)
        );

reg   lut_874_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_874_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_874_ff <= lut_874_out;
    end
end

assign out_data[874] = lut_874_ff;




// LUT : 875

wire lut_875_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101011111110000100001110001011010100111111000010001011011100),
            .DEVICE(DEVICE)
        )
    i_lut_875
        (
            .in_data({
                         in_data[384],
                         in_data[239],
                         in_data[773],
                         in_data[511],
                         in_data[375],
                         in_data[379]
                    }),
            .out_data(lut_875_out)
        );

reg   lut_875_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_875_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_875_ff <= lut_875_out;
    end
end

assign out_data[875] = lut_875_ff;




// LUT : 876

wire lut_876_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001100110111010010100001111101111011001111100111000100100100),
            .DEVICE(DEVICE)
        )
    i_lut_876
        (
            .in_data({
                         in_data[43],
                         in_data[586],
                         in_data[424],
                         in_data[209],
                         in_data[32],
                         in_data[104]
                    }),
            .out_data(lut_876_out)
        );

reg   lut_876_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_876_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_876_ff <= lut_876_out;
    end
end

assign out_data[876] = lut_876_ff;




// LUT : 877

wire lut_877_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010001110100101111110011100101011011111001001101000101011001),
            .DEVICE(DEVICE)
        )
    i_lut_877
        (
            .in_data({
                         in_data[169],
                         in_data[731],
                         in_data[203],
                         in_data[41],
                         in_data[21],
                         in_data[585]
                    }),
            .out_data(lut_877_out)
        );

reg   lut_877_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_877_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_877_ff <= lut_877_out;
    end
end

assign out_data[877] = lut_877_ff;




// LUT : 878

wire lut_878_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001101111011101001001010000110101000000010011100101101010001000),
            .DEVICE(DEVICE)
        )
    i_lut_878
        (
            .in_data({
                         in_data[198],
                         in_data[458],
                         in_data[38],
                         in_data[278],
                         in_data[436],
                         in_data[692]
                    }),
            .out_data(lut_878_out)
        );

reg   lut_878_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_878_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_878_ff <= lut_878_out;
    end
end

assign out_data[878] = lut_878_ff;




// LUT : 879

wire lut_879_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111010111111011011010011111100100011101110111010100100001011),
            .DEVICE(DEVICE)
        )
    i_lut_879
        (
            .in_data({
                         in_data[368],
                         in_data[284],
                         in_data[505],
                         in_data[470],
                         in_data[553],
                         in_data[776]
                    }),
            .out_data(lut_879_out)
        );

reg   lut_879_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_879_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_879_ff <= lut_879_out;
    end
end

assign out_data[879] = lut_879_ff;




// LUT : 880

wire lut_880_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000111111111000010010000111111111111111110100111101011111010),
            .DEVICE(DEVICE)
        )
    i_lut_880
        (
            .in_data({
                         in_data[70],
                         in_data[606],
                         in_data[249],
                         in_data[241],
                         in_data[343],
                         in_data[157]
                    }),
            .out_data(lut_880_out)
        );

reg   lut_880_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_880_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_880_ff <= lut_880_out;
    end
end

assign out_data[880] = lut_880_ff;




// LUT : 881

wire lut_881_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010111010111101110101111010100011010111110100010001000110101),
            .DEVICE(DEVICE)
        )
    i_lut_881
        (
            .in_data({
                         in_data[519],
                         in_data[777],
                         in_data[396],
                         in_data[409],
                         in_data[580],
                         in_data[374]
                    }),
            .out_data(lut_881_out)
        );

reg   lut_881_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_881_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_881_ff <= lut_881_out;
    end
end

assign out_data[881] = lut_881_ff;




// LUT : 882

wire lut_882_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001011011110100100110110110001101111100111010100101100010010000),
            .DEVICE(DEVICE)
        )
    i_lut_882
        (
            .in_data({
                         in_data[742],
                         in_data[108],
                         in_data[422],
                         in_data[6],
                         in_data[99],
                         in_data[72]
                    }),
            .out_data(lut_882_out)
        );

reg   lut_882_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_882_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_882_ff <= lut_882_out;
    end
end

assign out_data[882] = lut_882_ff;




// LUT : 883

wire lut_883_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110101011011001000000010001010101010011110110001001101110000),
            .DEVICE(DEVICE)
        )
    i_lut_883
        (
            .in_data({
                         in_data[80],
                         in_data[258],
                         in_data[119],
                         in_data[527],
                         in_data[383],
                         in_data[450]
                    }),
            .out_data(lut_883_out)
        );

reg   lut_883_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_883_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_883_ff <= lut_883_out;
    end
end

assign out_data[883] = lut_883_ff;




// LUT : 884

wire lut_884_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111010111111111110101011111111111111111111111100110000),
            .DEVICE(DEVICE)
        )
    i_lut_884
        (
            .in_data({
                         in_data[577],
                         in_data[576],
                         in_data[575],
                         in_data[548],
                         in_data[271],
                         in_data[600]
                    }),
            .out_data(lut_884_out)
        );

reg   lut_884_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_884_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_884_ff <= lut_884_out;
    end
end

assign out_data[884] = lut_884_ff;




// LUT : 885

wire lut_885_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011110001011110011011010100100001000000010111101011110101000),
            .DEVICE(DEVICE)
        )
    i_lut_885
        (
            .in_data({
                         in_data[659],
                         in_data[176],
                         in_data[48],
                         in_data[514],
                         in_data[517],
                         in_data[167]
                    }),
            .out_data(lut_885_out)
        );

reg   lut_885_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_885_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_885_ff <= lut_885_out;
    end
end

assign out_data[885] = lut_885_ff;




// LUT : 886

wire lut_886_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110111001000110111110001100101011101100001100101010110101110),
            .DEVICE(DEVICE)
        )
    i_lut_886
        (
            .in_data({
                         in_data[162],
                         in_data[555],
                         in_data[679],
                         in_data[582],
                         in_data[500],
                         in_data[0]
                    }),
            .out_data(lut_886_out)
        );

reg   lut_886_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_886_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_886_ff <= lut_886_out;
    end
end

assign out_data[886] = lut_886_ff;




// LUT : 887

wire lut_887_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011011010111110010011000100101010110000111011001010111011011),
            .DEVICE(DEVICE)
        )
    i_lut_887
        (
            .in_data({
                         in_data[55],
                         in_data[768],
                         in_data[559],
                         in_data[142],
                         in_data[488],
                         in_data[79]
                    }),
            .out_data(lut_887_out)
        );

reg   lut_887_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_887_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_887_ff <= lut_887_out;
    end
end

assign out_data[887] = lut_887_ff;




// LUT : 888

wire lut_888_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110001010110110100111010101101011000100110010001001001111111111),
            .DEVICE(DEVICE)
        )
    i_lut_888
        (
            .in_data({
                         in_data[378],
                         in_data[31],
                         in_data[344],
                         in_data[46],
                         in_data[10],
                         in_data[307]
                    }),
            .out_data(lut_888_out)
        );

reg   lut_888_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_888_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_888_ff <= lut_888_out;
    end
end

assign out_data[888] = lut_888_ff;




// LUT : 889

wire lut_889_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000011110101101101001111011100110011101010101011100100110000),
            .DEVICE(DEVICE)
        )
    i_lut_889
        (
            .in_data({
                         in_data[672],
                         in_data[225],
                         in_data[60],
                         in_data[2],
                         in_data[274],
                         in_data[570]
                    }),
            .out_data(lut_889_out)
        );

reg   lut_889_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_889_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_889_ff <= lut_889_out;
    end
end

assign out_data[889] = lut_889_ff;




// LUT : 890

wire lut_890_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101010100010001000001010100000001010100000001011001110111010),
            .DEVICE(DEVICE)
        )
    i_lut_890
        (
            .in_data({
                         in_data[668],
                         in_data[163],
                         in_data[318],
                         in_data[326],
                         in_data[211],
                         in_data[392]
                    }),
            .out_data(lut_890_out)
        );

reg   lut_890_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_890_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_890_ff <= lut_890_out;
    end
end

assign out_data[890] = lut_890_ff;




// LUT : 891

wire lut_891_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010110001111001010100110110101010101100001101010110100010100),
            .DEVICE(DEVICE)
        )
    i_lut_891
        (
            .in_data({
                         in_data[704],
                         in_data[110],
                         in_data[495],
                         in_data[633],
                         in_data[260],
                         in_data[448]
                    }),
            .out_data(lut_891_out)
        );

reg   lut_891_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_891_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_891_ff <= lut_891_out;
    end
end

assign out_data[891] = lut_891_ff;




// LUT : 892

wire lut_892_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000111001011111011110001100010011001001010100001000010101010),
            .DEVICE(DEVICE)
        )
    i_lut_892
        (
            .in_data({
                         in_data[377],
                         in_data[200],
                         in_data[332],
                         in_data[738],
                         in_data[547],
                         in_data[498]
                    }),
            .out_data(lut_892_out)
        );

reg   lut_892_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_892_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_892_ff <= lut_892_out;
    end
end

assign out_data[892] = lut_892_ff;




// LUT : 893

wire lut_893_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010101110000100010110010111100010110111111111001000110110111),
            .DEVICE(DEVICE)
        )
    i_lut_893
        (
            .in_data({
                         in_data[552],
                         in_data[336],
                         in_data[34],
                         in_data[116],
                         in_data[658],
                         in_data[607]
                    }),
            .out_data(lut_893_out)
        );

reg   lut_893_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_893_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_893_ff <= lut_893_out;
    end
end

assign out_data[893] = lut_893_ff;




// LUT : 894

wire lut_894_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001101011111100010011110101010110000010000000000101001110010100),
            .DEVICE(DEVICE)
        )
    i_lut_894
        (
            .in_data({
                         in_data[346],
                         in_data[172],
                         in_data[420],
                         in_data[574],
                         in_data[700],
                         in_data[740]
                    }),
            .out_data(lut_894_out)
        );

reg   lut_894_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_894_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_894_ff <= lut_894_out;
    end
end

assign out_data[894] = lut_894_ff;




// LUT : 895

wire lut_895_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011011010101111010100000001011011100011101110100111000110000),
            .DEVICE(DEVICE)
        )
    i_lut_895
        (
            .in_data({
                         in_data[432],
                         in_data[444],
                         in_data[131],
                         in_data[100],
                         in_data[454],
                         in_data[220]
                    }),
            .out_data(lut_895_out)
        );

reg   lut_895_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_895_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_895_ff <= lut_895_out;
    end
end

assign out_data[895] = lut_895_ff;




// LUT : 896

wire lut_896_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100011011100011010100011011010110010000000000000011101001011),
            .DEVICE(DEVICE)
        )
    i_lut_896
        (
            .in_data({
                         in_data[732],
                         in_data[733],
                         in_data[463],
                         in_data[75],
                         in_data[419],
                         in_data[402]
                    }),
            .out_data(lut_896_out)
        );

reg   lut_896_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_896_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_896_ff <= lut_896_out;
    end
end

assign out_data[896] = lut_896_ff;




// LUT : 897

wire lut_897_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011101000000111100111010100110010000010100110001110101010000000),
            .DEVICE(DEVICE)
        )
    i_lut_897
        (
            .in_data({
                         in_data[333],
                         in_data[12],
                         in_data[481],
                         in_data[88],
                         in_data[617],
                         in_data[604]
                    }),
            .out_data(lut_897_out)
        );

reg   lut_897_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_897_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_897_ff <= lut_897_out;
    end
end

assign out_data[897] = lut_897_ff;




// LUT : 898

wire lut_898_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111010100101001110110111011111111111111101110000011110010001),
            .DEVICE(DEVICE)
        )
    i_lut_898
        (
            .in_data({
                         in_data[416],
                         in_data[338],
                         in_data[287],
                         in_data[345],
                         in_data[350],
                         in_data[691]
                    }),
            .out_data(lut_898_out)
        );

reg   lut_898_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_898_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_898_ff <= lut_898_out;
    end
end

assign out_data[898] = lut_898_ff;




// LUT : 899

wire lut_899_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111010011001110000100111111111111011010011000011101111101111),
            .DEVICE(DEVICE)
        )
    i_lut_899
        (
            .in_data({
                         in_data[702],
                         in_data[188],
                         in_data[707],
                         in_data[597],
                         in_data[367],
                         in_data[173]
                    }),
            .out_data(lut_899_out)
        );

reg   lut_899_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_899_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_899_ff <= lut_899_out;
    end
end

assign out_data[899] = lut_899_ff;




// LUT : 900

wire lut_900_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111110001010100101000010011100010000000000000001000001001000001),
            .DEVICE(DEVICE)
        )
    i_lut_900
        (
            .in_data({
                         in_data[5],
                         in_data[496],
                         in_data[122],
                         in_data[558],
                         in_data[566],
                         in_data[536]
                    }),
            .out_data(lut_900_out)
        );

reg   lut_900_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_900_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_900_ff <= lut_900_out;
    end
end

assign out_data[900] = lut_900_ff;




// LUT : 901

wire lut_901_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111111001010000101010001111101001111111111110000111101001110),
            .DEVICE(DEVICE)
        )
    i_lut_901
        (
            .in_data({
                         in_data[710],
                         in_data[508],
                         in_data[373],
                         in_data[497],
                         in_data[236],
                         in_data[356]
                    }),
            .out_data(lut_901_out)
        );

reg   lut_901_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_901_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_901_ff <= lut_901_out;
    end
end

assign out_data[901] = lut_901_ff;




// LUT : 902

wire lut_902_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000101110010010110000101101000001101011011001101000101110101),
            .DEVICE(DEVICE)
        )
    i_lut_902
        (
            .in_data({
                         in_data[174],
                         in_data[65],
                         in_data[59],
                         in_data[723],
                         in_data[406],
                         in_data[22]
                    }),
            .out_data(lut_902_out)
        );

reg   lut_902_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_902_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_902_ff <= lut_902_out;
    end
end

assign out_data[902] = lut_902_ff;




// LUT : 903

wire lut_903_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101000111111000001001111010110111101001000111110110010100111),
            .DEVICE(DEVICE)
        )
    i_lut_903
        (
            .in_data({
                         in_data[299],
                         in_data[337],
                         in_data[696],
                         in_data[224],
                         in_data[47],
                         in_data[362]
                    }),
            .out_data(lut_903_out)
        );

reg   lut_903_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_903_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_903_ff <= lut_903_out;
    end
end

assign out_data[903] = lut_903_ff;




// LUT : 904

wire lut_904_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001111010011110101111001001101010100010011000100001101011100),
            .DEVICE(DEVICE)
        )
    i_lut_904
        (
            .in_data({
                         in_data[335],
                         in_data[369],
                         in_data[473],
                         in_data[613],
                         in_data[193],
                         in_data[764]
                    }),
            .out_data(lut_904_out)
        );

reg   lut_904_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_904_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_904_ff <= lut_904_out;
    end
end

assign out_data[904] = lut_904_ff;




// LUT : 905

wire lut_905_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010100001101000101010011010111010000110101010011011100110101),
            .DEVICE(DEVICE)
        )
    i_lut_905
        (
            .in_data({
                         in_data[195],
                         in_data[669],
                         in_data[665],
                         in_data[636],
                         in_data[265],
                         in_data[319]
                    }),
            .out_data(lut_905_out)
        );

reg   lut_905_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_905_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_905_ff <= lut_905_out;
    end
end

assign out_data[905] = lut_905_ff;




// LUT : 906

wire lut_906_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010101101001111000100110111000011011110011110000101100101111),
            .DEVICE(DEVICE)
        )
    i_lut_906
        (
            .in_data({
                         in_data[453],
                         in_data[645],
                         in_data[446],
                         in_data[471],
                         in_data[534],
                         in_data[50]
                    }),
            .out_data(lut_906_out)
        );

reg   lut_906_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_906_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_906_ff <= lut_906_out;
    end
end

assign out_data[906] = lut_906_ff;




// LUT : 907

wire lut_907_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010111001111010111010110111110000011101111010110001101101111),
            .DEVICE(DEVICE)
        )
    i_lut_907
        (
            .in_data({
                         in_data[73],
                         in_data[320],
                         in_data[61],
                         in_data[395],
                         in_data[708],
                         in_data[405]
                    }),
            .out_data(lut_907_out)
        );

reg   lut_907_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_907_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_907_ff <= lut_907_out;
    end
end

assign out_data[907] = lut_907_ff;




// LUT : 908

wire lut_908_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100101010110011101110001111010000010101101101100111111111110),
            .DEVICE(DEVICE)
        )
    i_lut_908
        (
            .in_data({
                         in_data[701],
                         in_data[515],
                         in_data[624],
                         in_data[58],
                         in_data[83],
                         in_data[151]
                    }),
            .out_data(lut_908_out)
        );

reg   lut_908_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_908_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_908_ff <= lut_908_out;
    end
end

assign out_data[908] = lut_908_ff;




// LUT : 909

wire lut_909_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001001110001000101111111110011110100011100100111011011111100),
            .DEVICE(DEVICE)
        )
    i_lut_909
        (
            .in_data({
                         in_data[538],
                         in_data[44],
                         in_data[729],
                         in_data[330],
                         in_data[366],
                         in_data[690]
                    }),
            .out_data(lut_909_out)
        );

reg   lut_909_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_909_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_909_ff <= lut_909_out;
    end
end

assign out_data[909] = lut_909_ff;




// LUT : 910

wire lut_910_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000011001000010011001100111111000101100010001000110011001111),
            .DEVICE(DEVICE)
        )
    i_lut_910
        (
            .in_data({
                         in_data[119],
                         in_data[383],
                         in_data[143],
                         in_data[465],
                         in_data[389],
                         in_data[118]
                    }),
            .out_data(lut_910_out)
        );

reg   lut_910_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_910_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_910_ff <= lut_910_out;
    end
end

assign out_data[910] = lut_910_ff;




// LUT : 911

wire lut_911_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101001000000010001001111001000001000000000000000001111111100001),
            .DEVICE(DEVICE)
        )
    i_lut_911
        (
            .in_data({
                         in_data[571],
                         in_data[152],
                         in_data[490],
                         in_data[477],
                         in_data[599],
                         in_data[754]
                    }),
            .out_data(lut_911_out)
        );

reg   lut_911_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_911_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_911_ff <= lut_911_out;
    end
end

assign out_data[911] = lut_911_ff;




// LUT : 912

wire lut_912_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111011111001100110000001100010110010010111111010001000010001),
            .DEVICE(DEVICE)
        )
    i_lut_912
        (
            .in_data({
                         in_data[429],
                         in_data[694],
                         in_data[398],
                         in_data[377],
                         in_data[43],
                         in_data[586]
                    }),
            .out_data(lut_912_out)
        );

reg   lut_912_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_912_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_912_ff <= lut_912_out;
    end
end

assign out_data[912] = lut_912_ff;




// LUT : 913

wire lut_913_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010110001001101100101010110011100110101111000011111000100101111),
            .DEVICE(DEVICE)
        )
    i_lut_913
        (
            .in_data({
                         in_data[67],
                         in_data[581],
                         in_data[716],
                         in_data[764],
                         in_data[86],
                         in_data[216]
                    }),
            .out_data(lut_913_out)
        );

reg   lut_913_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_913_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_913_ff <= lut_913_out;
    end
end

assign out_data[913] = lut_913_ff;




// LUT : 914

wire lut_914_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000110001010101111000111001011001000011000111101110000011001),
            .DEVICE(DEVICE)
        )
    i_lut_914
        (
            .in_data({
                         in_data[706],
                         in_data[664],
                         in_data[592],
                         in_data[54],
                         in_data[558],
                         in_data[507]
                    }),
            .out_data(lut_914_out)
        );

reg   lut_914_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_914_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_914_ff <= lut_914_out;
    end
end

assign out_data[914] = lut_914_ff;




// LUT : 915

wire lut_915_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010011010000101011100110001000011010001010100010001100010010),
            .DEVICE(DEVICE)
        )
    i_lut_915
        (
            .in_data({
                         in_data[193],
                         in_data[76],
                         in_data[608],
                         in_data[302],
                         in_data[122],
                         in_data[451]
                    }),
            .out_data(lut_915_out)
        );

reg   lut_915_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_915_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_915_ff <= lut_915_out;
    end
end

assign out_data[915] = lut_915_ff;




// LUT : 916

wire lut_916_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100101001111011001011110110001010101011101100011100111000001010),
            .DEVICE(DEVICE)
        )
    i_lut_916
        (
            .in_data({
                         in_data[425],
                         in_data[26],
                         in_data[501],
                         in_data[205],
                         in_data[336],
                         in_data[357]
                    }),
            .out_data(lut_916_out)
        );

reg   lut_916_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_916_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_916_ff <= lut_916_out;
    end
end

assign out_data[916] = lut_916_ff;




// LUT : 917

wire lut_917_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000110100011111100100101001010100000000000001011000001000000),
            .DEVICE(DEVICE)
        )
    i_lut_917
        (
            .in_data({
                         in_data[483],
                         in_data[346],
                         in_data[153],
                         in_data[63],
                         in_data[330],
                         in_data[433]
                    }),
            .out_data(lut_917_out)
        );

reg   lut_917_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_917_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_917_ff <= lut_917_out;
    end
end

assign out_data[917] = lut_917_ff;




// LUT : 918

wire lut_918_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100101110110010000001000100111011001101101100010110010111011),
            .DEVICE(DEVICE)
        )
    i_lut_918
        (
            .in_data({
                         in_data[709],
                         in_data[280],
                         in_data[566],
                         in_data[715],
                         in_data[222],
                         in_data[141]
                    }),
            .out_data(lut_918_out)
        );

reg   lut_918_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_918_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_918_ff <= lut_918_out;
    end
end

assign out_data[918] = lut_918_ff;




// LUT : 919

wire lut_919_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000011010110111111011100000011010011000000001001110000101000011),
            .DEVICE(DEVICE)
        )
    i_lut_919
        (
            .in_data({
                         in_data[130],
                         in_data[172],
                         in_data[375],
                         in_data[278],
                         in_data[40],
                         in_data[611]
                    }),
            .out_data(lut_919_out)
        );

reg   lut_919_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_919_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_919_ff <= lut_919_out;
    end
end

assign out_data[919] = lut_919_ff;




// LUT : 920

wire lut_920_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110011101110010011100000010111100101000000010001100101110100011),
            .DEVICE(DEVICE)
        )
    i_lut_920
        (
            .in_data({
                         in_data[618],
                         in_data[292],
                         in_data[755],
                         in_data[583],
                         in_data[369],
                         in_data[604]
                    }),
            .out_data(lut_920_out)
        );

reg   lut_920_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_920_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_920_ff <= lut_920_out;
    end
end

assign out_data[920] = lut_920_ff;




// LUT : 921

wire lut_921_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001100110111111101110010111001010111001000111110010000010100000),
            .DEVICE(DEVICE)
        )
    i_lut_921
        (
            .in_data({
                         in_data[531],
                         in_data[352],
                         in_data[394],
                         in_data[349],
                         in_data[609],
                         in_data[728]
                    }),
            .out_data(lut_921_out)
        );

reg   lut_921_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_921_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_921_ff <= lut_921_out;
    end
end

assign out_data[921] = lut_921_ff;




// LUT : 922

wire lut_922_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100111110101011001101111101011100010011000000001110110000100),
            .DEVICE(DEVICE)
        )
    i_lut_922
        (
            .in_data({
                         in_data[17],
                         in_data[712],
                         in_data[475],
                         in_data[347],
                         in_data[89],
                         in_data[70]
                    }),
            .out_data(lut_922_out)
        );

reg   lut_922_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_922_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_922_ff <= lut_922_out;
    end
end

assign out_data[922] = lut_922_ff;




// LUT : 923

wire lut_923_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000111100101000001100000101011010100011101100111101001101010),
            .DEVICE(DEVICE)
        )
    i_lut_923
        (
            .in_data({
                         in_data[550],
                         in_data[700],
                         in_data[750],
                         in_data[214],
                         in_data[773],
                         in_data[27]
                    }),
            .out_data(lut_923_out)
        );

reg   lut_923_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_923_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_923_ff <= lut_923_out;
    end
end

assign out_data[923] = lut_923_ff;




// LUT : 924

wire lut_924_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111001010010000101010111100101001000000010001100111111001001),
            .DEVICE(DEVICE)
        )
    i_lut_924
        (
            .in_data({
                         in_data[617],
                         in_data[179],
                         in_data[406],
                         in_data[530],
                         in_data[331],
                         in_data[326]
                    }),
            .out_data(lut_924_out)
        );

reg   lut_924_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_924_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_924_ff <= lut_924_out;
    end
end

assign out_data[924] = lut_924_ff;




// LUT : 925

wire lut_925_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101111110100111001000001100111011010001010001111001000101000),
            .DEVICE(DEVICE)
        )
    i_lut_925
        (
            .in_data({
                         in_data[536],
                         in_data[38],
                         in_data[224],
                         in_data[461],
                         in_data[460],
                         in_data[195]
                    }),
            .out_data(lut_925_out)
        );

reg   lut_925_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_925_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_925_ff <= lut_925_out;
    end
end

assign out_data[925] = lut_925_ff;




// LUT : 926

wire lut_926_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111101000011101111100110111001000011100111101001010001110000),
            .DEVICE(DEVICE)
        )
    i_lut_926
        (
            .in_data({
                         in_data[509],
                         in_data[420],
                         in_data[177],
                         in_data[484],
                         in_data[225],
                         in_data[693]
                    }),
            .out_data(lut_926_out)
        );

reg   lut_926_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_926_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_926_ff <= lut_926_out;
    end
end

assign out_data[926] = lut_926_ff;




// LUT : 927

wire lut_927_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100101100010111001001110101010110110101010010100011100100110110),
            .DEVICE(DEVICE)
        )
    i_lut_927
        (
            .in_data({
                         in_data[680],
                         in_data[11],
                         in_data[229],
                         in_data[668],
                         in_data[50],
                         in_data[64]
                    }),
            .out_data(lut_927_out)
        );

reg   lut_927_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_927_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_927_ff <= lut_927_out;
    end
end

assign out_data[927] = lut_927_ff;




// LUT : 928

wire lut_928_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010001001111111100111110010010100001101010110101000011011101),
            .DEVICE(DEVICE)
        )
    i_lut_928
        (
            .in_data({
                         in_data[206],
                         in_data[370],
                         in_data[707],
                         in_data[691],
                         in_data[714],
                         in_data[576]
                    }),
            .out_data(lut_928_out)
        );

reg   lut_928_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_928_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_928_ff <= lut_928_out;
    end
end

assign out_data[928] = lut_928_ff;




// LUT : 929

wire lut_929_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001011101100011101011111011101011111000000001100111000001111),
            .DEVICE(DEVICE)
        )
    i_lut_929
        (
            .in_data({
                         in_data[434],
                         in_data[685],
                         in_data[758],
                         in_data[293],
                         in_data[316],
                         in_data[464]
                    }),
            .out_data(lut_929_out)
        );

reg   lut_929_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_929_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_929_ff <= lut_929_out;
    end
end

assign out_data[929] = lut_929_ff;




// LUT : 930

wire lut_930_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000110101001110101011001111011011011011110100001111111011010000),
            .DEVICE(DEVICE)
        )
    i_lut_930
        (
            .in_data({
                         in_data[512],
                         in_data[84],
                         in_data[323],
                         in_data[546],
                         in_data[516],
                         in_data[81]
                    }),
            .out_data(lut_930_out)
        );

reg   lut_930_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_930_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_930_ff <= lut_930_out;
    end
end

assign out_data[930] = lut_930_ff;




// LUT : 931

wire lut_931_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001010010000100110101100100010001000100000010000100010100001),
            .DEVICE(DEVICE)
        )
    i_lut_931
        (
            .in_data({
                         in_data[564],
                         in_data[208],
                         in_data[178],
                         in_data[47],
                         in_data[129],
                         in_data[80]
                    }),
            .out_data(lut_931_out)
        );

reg   lut_931_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_931_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_931_ff <= lut_931_out;
    end
end

assign out_data[931] = lut_931_ff;




// LUT : 932

wire lut_932_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110011000001011100011110111000010100010000000111100001001000011),
            .DEVICE(DEVICE)
        )
    i_lut_932
        (
            .in_data({
                         in_data[159],
                         in_data[652],
                         in_data[110],
                         in_data[743],
                         in_data[97],
                         in_data[413]
                    }),
            .out_data(lut_932_out)
        );

reg   lut_932_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_932_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_932_ff <= lut_932_out;
    end
end

assign out_data[932] = lut_932_ff;




// LUT : 933

wire lut_933_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010111100100011000000011011001111101011010000100011111010111110),
            .DEVICE(DEVICE)
        )
    i_lut_933
        (
            .in_data({
                         in_data[747],
                         in_data[757],
                         in_data[416],
                         in_data[21],
                         in_data[527],
                         in_data[543]
                    }),
            .out_data(lut_933_out)
        );

reg   lut_933_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_933_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_933_ff <= lut_933_out;
    end
end

assign out_data[933] = lut_933_ff;




// LUT : 934

wire lut_934_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111100011100100110111000011010001101010010001100011001011010110),
            .DEVICE(DEVICE)
        )
    i_lut_934
        (
            .in_data({
                         in_data[22],
                         in_data[262],
                         in_data[596],
                         in_data[468],
                         in_data[740],
                         in_data[724]
                    }),
            .out_data(lut_934_out)
        );

reg   lut_934_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_934_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_934_ff <= lut_934_out;
    end
end

assign out_data[934] = lut_934_ff;




// LUT : 935

wire lut_935_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011101000100101101000111110001110001011100101110111000111011010),
            .DEVICE(DEVICE)
        )
    i_lut_935
        (
            .in_data({
                         in_data[82],
                         in_data[244],
                         in_data[616],
                         in_data[339],
                         in_data[414],
                         in_data[649]
                    }),
            .out_data(lut_935_out)
        );

reg   lut_935_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_935_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_935_ff <= lut_935_out;
    end
end

assign out_data[935] = lut_935_ff;




// LUT : 936

wire lut_936_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000010111110111111001100101011010010001011110101100000101011),
            .DEVICE(DEVICE)
        )
    i_lut_936
        (
            .in_data({
                         in_data[215],
                         in_data[299],
                         in_data[335],
                         in_data[761],
                         in_data[573],
                         in_data[521]
                    }),
            .out_data(lut_936_out)
        );

reg   lut_936_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_936_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_936_ff <= lut_936_out;
    end
end

assign out_data[936] = lut_936_ff;




// LUT : 937

wire lut_937_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011110011111000011110000010000101111000011000001111000100100),
            .DEVICE(DEVICE)
        )
    i_lut_937
        (
            .in_data({
                         in_data[241],
                         in_data[582],
                         in_data[517],
                         in_data[478],
                         in_data[600],
                         in_data[212]
                    }),
            .out_data(lut_937_out)
        );

reg   lut_937_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_937_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_937_ff <= lut_937_out;
    end
end

assign out_data[937] = lut_937_ff;




// LUT : 938

wire lut_938_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101010010101100111101101110100111010100101011111010110011000),
            .DEVICE(DEVICE)
        )
    i_lut_938
        (
            .in_data({
                         in_data[471],
                         in_data[271],
                         in_data[480],
                         in_data[486],
                         in_data[113],
                         in_data[145]
                    }),
            .out_data(lut_938_out)
        );

reg   lut_938_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_938_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_938_ff <= lut_938_out;
    end
end

assign out_data[938] = lut_938_ff;




// LUT : 939

wire lut_939_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101100101010001100011011100101110110011101110000001000110011010),
            .DEVICE(DEVICE)
        )
    i_lut_939
        (
            .in_data({
                         in_data[197],
                         in_data[380],
                         in_data[771],
                         in_data[458],
                         in_data[646],
                         in_data[16]
                    }),
            .out_data(lut_939_out)
        );

reg   lut_939_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_939_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_939_ff <= lut_939_out;
    end
end

assign out_data[939] = lut_939_ff;




// LUT : 940

wire lut_940_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001110000001110110001010001011101001000101100000111111001001111),
            .DEVICE(DEVICE)
        )
    i_lut_940
        (
            .in_data({
                         in_data[114],
                         in_data[588],
                         in_data[345],
                         in_data[777],
                         in_data[597],
                         in_data[137]
                    }),
            .out_data(lut_940_out)
        );

reg   lut_940_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_940_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_940_ff <= lut_940_out;
    end
end

assign out_data[940] = lut_940_ff;




// LUT : 941

wire lut_941_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110110000000000100100001100010111010000010000011101000000000101),
            .DEVICE(DEVICE)
        )
    i_lut_941
        (
            .in_data({
                         in_data[628],
                         in_data[542],
                         in_data[147],
                         in_data[447],
                         in_data[631],
                         in_data[228]
                    }),
            .out_data(lut_941_out)
        );

reg   lut_941_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_941_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_941_ff <= lut_941_out;
    end
end

assign out_data[941] = lut_941_ff;




// LUT : 942

wire lut_942_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111100011110000011111001111100111011111110001110111101101100),
            .DEVICE(DEVICE)
        )
    i_lut_942
        (
            .in_data({
                         in_data[73],
                         in_data[683],
                         in_data[259],
                         in_data[312],
                         in_data[117],
                         in_data[630]
                    }),
            .out_data(lut_942_out)
        );

reg   lut_942_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_942_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_942_ff <= lut_942_out;
    end
end

assign out_data[942] = lut_942_ff;




// LUT : 943

wire lut_943_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110110010001001101010000111111101000100110110111000001000100),
            .DEVICE(DEVICE)
        )
    i_lut_943
        (
            .in_data({
                         in_data[538],
                         in_data[282],
                         in_data[182],
                         in_data[340],
                         in_data[696],
                         in_data[602]
                    }),
            .out_data(lut_943_out)
        );

reg   lut_943_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_943_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_943_ff <= lut_943_out;
    end
end

assign out_data[943] = lut_943_ff;




// LUT : 944

wire lut_944_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101001011000001010101001100000000100010000001110100110110001),
            .DEVICE(DEVICE)
        )
    i_lut_944
        (
            .in_data({
                         in_data[171],
                         in_data[635],
                         in_data[595],
                         in_data[660],
                         in_data[614],
                         in_data[92]
                    }),
            .out_data(lut_944_out)
        );

reg   lut_944_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_944_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_944_ff <= lut_944_out;
    end
end

assign out_data[944] = lut_944_ff;




// LUT : 945

wire lut_945_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000111111011100111011101111111011011000111111011011010011111),
            .DEVICE(DEVICE)
        )
    i_lut_945
        (
            .in_data({
                         in_data[513],
                         in_data[496],
                         in_data[237],
                         in_data[277],
                         in_data[18],
                         in_data[7]
                    }),
            .out_data(lut_945_out)
        );

reg   lut_945_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_945_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_945_ff <= lut_945_out;
    end
end

assign out_data[945] = lut_945_ff;




// LUT : 946

wire lut_946_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010110001011010111111001010000001001000001110100111111100011111),
            .DEVICE(DEVICE)
        )
    i_lut_946
        (
            .in_data({
                         in_data[128],
                         in_data[367],
                         in_data[372],
                         in_data[734],
                         in_data[246],
                         in_data[65]
                    }),
            .out_data(lut_946_out)
        );

reg   lut_946_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_946_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_946_ff <= lut_946_out;
    end
end

assign out_data[946] = lut_946_ff;




// LUT : 947

wire lut_947_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000100011000000001000011011111101001001100011111110110111100),
            .DEVICE(DEVICE)
        )
    i_lut_947
        (
            .in_data({
                         in_data[120],
                         in_data[167],
                         in_data[165],
                         in_data[637],
                         in_data[624],
                         in_data[258]
                    }),
            .out_data(lut_947_out)
        );

reg   lut_947_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_947_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_947_ff <= lut_947_out;
    end
end

assign out_data[947] = lut_947_ff;




// LUT : 948

wire lut_948_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000000100110011101001000000001001101100010001000011001001011),
            .DEVICE(DEVICE)
        )
    i_lut_948
        (
            .in_data({
                         in_data[180],
                         in_data[226],
                         in_data[421],
                         in_data[284],
                         in_data[33],
                         in_data[679]
                    }),
            .out_data(lut_948_out)
        );

reg   lut_948_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_948_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_948_ff <= lut_948_out;
    end
end

assign out_data[948] = lut_948_ff;




// LUT : 949

wire lut_949_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111101011001110100110101100011100011001111110010011001110101),
            .DEVICE(DEVICE)
        )
    i_lut_949
        (
            .in_data({
                         in_data[391],
                         in_data[88],
                         in_data[762],
                         in_data[674],
                         in_data[437],
                         in_data[540]
                    }),
            .out_data(lut_949_out)
        );

reg   lut_949_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_949_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_949_ff <= lut_949_out;
    end
end

assign out_data[949] = lut_949_ff;




// LUT : 950

wire lut_950_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011100110010110110100011111111101110000010110000011110101010),
            .DEVICE(DEVICE)
        )
    i_lut_950
        (
            .in_data({
                         in_data[502],
                         in_data[650],
                         in_data[725],
                         in_data[470],
                         in_data[622],
                         in_data[102]
                    }),
            .out_data(lut_950_out)
        );

reg   lut_950_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_950_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_950_ff <= lut_950_out;
    end
end

assign out_data[950] = lut_950_ff;




// LUT : 951

wire lut_951_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100011101101100000011111001001011001100000010011100110001011011),
            .DEVICE(DEVICE)
        )
    i_lut_951
        (
            .in_data({
                         in_data[68],
                         in_data[231],
                         in_data[711],
                         in_data[654],
                         in_data[473],
                         in_data[663]
                    }),
            .out_data(lut_951_out)
        );

reg   lut_951_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_951_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_951_ff <= lut_951_out;
    end
end

assign out_data[951] = lut_951_ff;




// LUT : 952

wire lut_952_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110011101110100101011111101101011010110010101001101010000000100),
            .DEVICE(DEVICE)
        )
    i_lut_952
        (
            .in_data({
                         in_data[71],
                         in_data[603],
                         in_data[234],
                         in_data[121],
                         in_data[488],
                         in_data[390]
                    }),
            .out_data(lut_952_out)
        );

reg   lut_952_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_952_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_952_ff <= lut_952_out;
    end
end

assign out_data[952] = lut_952_ff;




// LUT : 953

wire lut_953_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010101000010111001110001100100011011111111010000101101011111),
            .DEVICE(DEVICE)
        )
    i_lut_953
        (
            .in_data({
                         in_data[642],
                         in_data[45],
                         in_data[242],
                         in_data[360],
                         in_data[733],
                         in_data[79]
                    }),
            .out_data(lut_953_out)
        );

reg   lut_953_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_953_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_953_ff <= lut_953_out;
    end
end

assign out_data[953] = lut_953_ff;




// LUT : 954

wire lut_954_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010100001100010011000100000010010000001000001111101001001010),
            .DEVICE(DEVICE)
        )
    i_lut_954
        (
            .in_data({
                         in_data[708],
                         in_data[769],
                         in_data[522],
                         in_data[499],
                         in_data[511],
                         in_data[457]
                    }),
            .out_data(lut_954_out)
        );

reg   lut_954_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_954_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_954_ff <= lut_954_out;
    end
end

assign out_data[954] = lut_954_ff;




// LUT : 955

wire lut_955_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111001000110110000001000010010101110100001000100100001000010),
            .DEVICE(DEVICE)
        )
    i_lut_955
        (
            .in_data({
                         in_data[199],
                         in_data[395],
                         in_data[767],
                         in_data[55],
                         in_data[574],
                         in_data[127]
                    }),
            .out_data(lut_955_out)
        );

reg   lut_955_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_955_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_955_ff <= lut_955_out;
    end
end

assign out_data[955] = lut_955_ff;




// LUT : 956

wire lut_956_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011001001111110010000111100100110111111101110100001011000110),
            .DEVICE(DEVICE)
        )
    i_lut_956
        (
            .in_data({
                         in_data[446],
                         in_data[131],
                         in_data[657],
                         in_data[396],
                         in_data[78],
                         in_data[90]
                    }),
            .out_data(lut_956_out)
        );

reg   lut_956_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_956_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_956_ff <= lut_956_out;
    end
end

assign out_data[956] = lut_956_ff;




// LUT : 957

wire lut_957_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001110011011100001000011101101010101001110011101011100000100),
            .DEVICE(DEVICE)
        )
    i_lut_957
        (
            .in_data({
                         in_data[772],
                         in_data[658],
                         in_data[686],
                         in_data[489],
                         in_data[621],
                         in_data[104]
                    }),
            .out_data(lut_957_out)
        );

reg   lut_957_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_957_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_957_ff <= lut_957_out;
    end
end

assign out_data[957] = lut_957_ff;




// LUT : 958

wire lut_958_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101101011101111001100100101000000000001111110010001000101110),
            .DEVICE(DEVICE)
        )
    i_lut_958
        (
            .in_data({
                         in_data[9],
                         in_data[682],
                         in_data[452],
                         in_data[426],
                         in_data[238],
                         in_data[322]
                    }),
            .out_data(lut_958_out)
        );

reg   lut_958_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_958_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_958_ff <= lut_958_out;
    end
end

assign out_data[958] = lut_958_ff;




// LUT : 959

wire lut_959_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011100111001000011011100000010101000001110110000111111111010),
            .DEVICE(DEVICE)
        )
    i_lut_959
        (
            .in_data({
                         in_data[405],
                         in_data[569],
                         in_data[3],
                         in_data[577],
                         in_data[732],
                         in_data[155]
                    }),
            .out_data(lut_959_out)
        );

reg   lut_959_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_959_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_959_ff <= lut_959_out;
    end
end

assign out_data[959] = lut_959_ff;




// LUT : 960

wire lut_960_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011100011111111110110011111000010000010011111111101111101110000),
            .DEVICE(DEVICE)
        )
    i_lut_960
        (
            .in_data({
                         in_data[350],
                         in_data[173],
                         in_data[387],
                         in_data[297],
                         in_data[181],
                         in_data[106]
                    }),
            .out_data(lut_960_out)
        );

reg   lut_960_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_960_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_960_ff <= lut_960_out;
    end
end

assign out_data[960] = lut_960_ff;




// LUT : 961

wire lut_961_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110100010101000111101001110010000100000101110111111010110110101),
            .DEVICE(DEVICE)
        )
    i_lut_961
        (
            .in_data({
                         in_data[93],
                         in_data[626],
                         in_data[427],
                         in_data[28],
                         in_data[697],
                         in_data[373]
                    }),
            .out_data(lut_961_out)
        );

reg   lut_961_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_961_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_961_ff <= lut_961_out;
    end
end

assign out_data[961] = lut_961_ff;




// LUT : 962

wire lut_962_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000011101101011001100101011111010101000101001101010111111000),
            .DEVICE(DEVICE)
        )
    i_lut_962
        (
            .in_data({
                         in_data[66],
                         in_data[25],
                         in_data[741],
                         in_data[296],
                         in_data[239],
                         in_data[5]
                    }),
            .out_data(lut_962_out)
        );

reg   lut_962_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_962_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_962_ff <= lut_962_out;
    end
end

assign out_data[962] = lut_962_ff;




// LUT : 963

wire lut_963_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000110110100000011100010010111010101101110011101001010111011100),
            .DEVICE(DEVICE)
        )
    i_lut_963
        (
            .in_data({
                         in_data[148],
                         in_data[412],
                         in_data[781],
                         in_data[525],
                         in_data[32],
                         in_data[307]
                    }),
            .out_data(lut_963_out)
        );

reg   lut_963_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_963_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_963_ff <= lut_963_out;
    end
end

assign out_data[963] = lut_963_ff;




// LUT : 964

wire lut_964_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100010100001100000000000000000110111001001100011000000010000001),
            .DEVICE(DEVICE)
        )
    i_lut_964
        (
            .in_data({
                         in_data[184],
                         in_data[532],
                         in_data[514],
                         in_data[72],
                         in_data[329],
                         in_data[612]
                    }),
            .out_data(lut_964_out)
        );

reg   lut_964_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_964_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_964_ff <= lut_964_out;
    end
end

assign out_data[964] = lut_964_ff;




// LUT : 965

wire lut_965_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110010100010010110101010010001101000110000000000000010100001001),
            .DEVICE(DEVICE)
        )
    i_lut_965
        (
            .in_data({
                         in_data[343],
                         in_data[607],
                         in_data[107],
                         in_data[176],
                         in_data[619],
                         in_data[146]
                    }),
            .out_data(lut_965_out)
        );

reg   lut_965_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_965_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_965_ff <= lut_965_out;
    end
end

assign out_data[965] = lut_965_ff;




// LUT : 966

wire lut_966_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111100101111010011111101111101101010000011111101011100010111),
            .DEVICE(DEVICE)
        )
    i_lut_966
        (
            .in_data({
                         in_data[435],
                         in_data[625],
                         in_data[485],
                         in_data[645],
                         in_data[469],
                         in_data[194]
                    }),
            .out_data(lut_966_out)
        );

reg   lut_966_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_966_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_966_ff <= lut_966_out;
    end
end

assign out_data[966] = lut_966_ff;




// LUT : 967

wire lut_967_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010101010111100001111001011100110111010001111000011111000000),
            .DEVICE(DEVICE)
        )
    i_lut_967
        (
            .in_data({
                         in_data[556],
                         in_data[472],
                         in_data[584],
                         in_data[319],
                         in_data[261],
                         in_data[96]
                    }),
            .out_data(lut_967_out)
        );

reg   lut_967_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_967_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_967_ff <= lut_967_out;
    end
end

assign out_data[967] = lut_967_ff;




// LUT : 968

wire lut_968_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001000111100010101010000001000100001110011110000101100101001),
            .DEVICE(DEVICE)
        )
    i_lut_968
        (
            .in_data({
                         in_data[589],
                         in_data[783],
                         in_data[166],
                         in_data[187],
                         in_data[424],
                         in_data[731]
                    }),
            .out_data(lut_968_out)
        );

reg   lut_968_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_968_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_968_ff <= lut_968_out;
    end
end

assign out_data[968] = lut_968_ff;




// LUT : 969

wire lut_969_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110010100000011111101111011011111101000111111110010111100000101),
            .DEVICE(DEVICE)
        )
    i_lut_969
        (
            .in_data({
                         in_data[776],
                         in_data[647],
                         in_data[570],
                         in_data[407],
                         in_data[467],
                         in_data[547]
                    }),
            .out_data(lut_969_out)
        );

reg   lut_969_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_969_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_969_ff <= lut_969_out;
    end
end

assign out_data[969] = lut_969_ff;




// LUT : 970

wire lut_970_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001010000101101110110010101111111010000110001001101111001111),
            .DEVICE(DEVICE)
        )
    i_lut_970
        (
            .in_data({
                         in_data[233],
                         in_data[132],
                         in_data[174],
                         in_data[0],
                         in_data[4],
                         in_data[219]
                    }),
            .out_data(lut_970_out)
        );

reg   lut_970_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_970_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_970_ff <= lut_970_out;
    end
end

assign out_data[970] = lut_970_ff;




// LUT : 971

wire lut_971_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111101111111111111111100110011111111011111111111111111001100),
            .DEVICE(DEVICE)
        )
    i_lut_971
        (
            .in_data({
                         in_data[431],
                         in_data[48],
                         in_data[440],
                         in_data[269],
                         in_data[382],
                         in_data[211]
                    }),
            .out_data(lut_971_out)
        );

reg   lut_971_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_971_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_971_ff <= lut_971_out;
    end
end

assign out_data[971] = lut_971_ff;




// LUT : 972

wire lut_972_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000000010000111100000001000010010000001100001101001011100011),
            .DEVICE(DEVICE)
        )
    i_lut_972
        (
            .in_data({
                         in_data[738],
                         in_data[710],
                         in_data[371],
                         in_data[20],
                         in_data[315],
                         in_data[213]
                    }),
            .out_data(lut_972_out)
        );

reg   lut_972_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_972_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_972_ff <= lut_972_out;
    end
end

assign out_data[972] = lut_972_ff;




// LUT : 973

wire lut_973_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100001001101011111111101100000101110011101111011010010111000),
            .DEVICE(DEVICE)
        )
    i_lut_973
        (
            .in_data({
                         in_data[644],
                         in_data[317],
                         in_data[295],
                         in_data[698],
                         in_data[53],
                         in_data[286]
                    }),
            .out_data(lut_973_out)
        );

reg   lut_973_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_973_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_973_ff <= lut_973_out;
    end
end

assign out_data[973] = lut_973_ff;




// LUT : 974

wire lut_974_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111001111110111111111001101010111110011100100111111100011111),
            .DEVICE(DEVICE)
        )
    i_lut_974
        (
            .in_data({
                         in_data[409],
                         in_data[419],
                         in_data[459],
                         in_data[669],
                         in_data[684],
                         in_data[585]
                    }),
            .out_data(lut_974_out)
        );

reg   lut_974_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_974_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_974_ff <= lut_974_out;
    end
end

assign out_data[974] = lut_974_ff;




// LUT : 975

wire lut_975_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010100101010011100100100101000100001011000001010000100100000),
            .DEVICE(DEVICE)
        )
    i_lut_975
        (
            .in_data({
                         in_data[775],
                         in_data[365],
                         in_data[359],
                         in_data[670],
                         in_data[423],
                         in_data[202]
                    }),
            .out_data(lut_975_out)
        );

reg   lut_975_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_975_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_975_ff <= lut_975_out;
    end
end

assign out_data[975] = lut_975_ff;




// LUT : 976

wire lut_976_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011100001111011011111101101001010000100011111000111110001000),
            .DEVICE(DEVICE)
        )
    i_lut_976
        (
            .in_data({
                         in_data[287],
                         in_data[341],
                         in_data[249],
                         in_data[112],
                         in_data[601],
                         in_data[388]
                    }),
            .out_data(lut_976_out)
        );

reg   lut_976_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_976_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_976_ff <= lut_976_out;
    end
end

assign out_data[976] = lut_976_ff;




// LUT : 977

wire lut_977_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101001111110101000101110101000000110010110111010101010100000),
            .DEVICE(DEVICE)
        )
    i_lut_977
        (
            .in_data({
                         in_data[492],
                         in_data[503],
                         in_data[411],
                         in_data[450],
                         in_data[34],
                         in_data[665]
                    }),
            .out_data(lut_977_out)
        );

reg   lut_977_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_977_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_977_ff <= lut_977_out;
    end
end

assign out_data[977] = lut_977_ff;




// LUT : 978

wire lut_978_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110101000010001011101110010011101100101101111111111111110101111),
            .DEVICE(DEVICE)
        )
    i_lut_978
        (
            .in_data({
                         in_data[268],
                         in_data[560],
                         in_data[313],
                         in_data[175],
                         in_data[661],
                         in_data[283]
                    }),
            .out_data(lut_978_out)
        );

reg   lut_978_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_978_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_978_ff <= lut_978_out;
    end
end

assign out_data[978] = lut_978_ff;




// LUT : 979

wire lut_979_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101010101010011110010100100111110010101101111111100001111000),
            .DEVICE(DEVICE)
        )
    i_lut_979
        (
            .in_data({
                         in_data[515],
                         in_data[636],
                         in_data[385],
                         in_data[578],
                         in_data[756],
                         in_data[91]
                    }),
            .out_data(lut_979_out)
        );

reg   lut_979_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_979_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_979_ff <= lut_979_out;
    end
end

assign out_data[979] = lut_979_ff;




// LUT : 980

wire lut_980_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110000000100101010111000111100001100000010000000000011011100),
            .DEVICE(DEVICE)
        )
    i_lut_980
        (
            .in_data({
                         in_data[403],
                         in_data[506],
                         in_data[217],
                         in_data[133],
                         in_data[162],
                         in_data[263]
                    }),
            .out_data(lut_980_out)
        );

reg   lut_980_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_980_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_980_ff <= lut_980_out;
    end
end

assign out_data[980] = lut_980_ff;




// LUT : 981

wire lut_981_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011100101001110110111101011000111111011101101101111001010010111),
            .DEVICE(DEVICE)
        )
    i_lut_981
        (
            .in_data({
                         in_data[487],
                         in_data[445],
                         in_data[157],
                         in_data[332],
                         in_data[753],
                         in_data[422]
                    }),
            .out_data(lut_981_out)
        );

reg   lut_981_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_981_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_981_ff <= lut_981_out;
    end
end

assign out_data[981] = lut_981_ff;




// LUT : 982

wire lut_982_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110011011010111111101000010100010111010101010110100010111111),
            .DEVICE(DEVICE)
        )
    i_lut_982
        (
            .in_data({
                         in_data[766],
                         in_data[46],
                         in_data[439],
                         in_data[415],
                         in_data[505],
                         in_data[30]
                    }),
            .out_data(lut_982_out)
        );

reg   lut_982_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_982_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_982_ff <= lut_982_out;
    end
end

assign out_data[982] = lut_982_ff;




// LUT : 983

wire lut_983_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111000001101000001110100010011111111011111110110111110001100),
            .DEVICE(DEVICE)
        )
    i_lut_983
        (
            .in_data({
                         in_data[565],
                         in_data[720],
                         in_data[526],
                         in_data[138],
                         in_data[554],
                         in_data[721]
                    }),
            .out_data(lut_983_out)
        );

reg   lut_983_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_983_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_983_ff <= lut_983_out;
    end
end

assign out_data[983] = lut_983_ff;




// LUT : 984

wire lut_984_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000000000000110101010010110001010001101100011111101010001010),
            .DEVICE(DEVICE)
        )
    i_lut_984
        (
            .in_data({
                         in_data[479],
                         in_data[35],
                         in_data[676],
                         in_data[311],
                         in_data[651],
                         in_data[404]
                    }),
            .out_data(lut_984_out)
        );

reg   lut_984_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_984_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_984_ff <= lut_984_out;
    end
end

assign out_data[984] = lut_984_ff;




// LUT : 985

wire lut_985_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000001110000001110000110100001101101110111101100111111110010),
            .DEVICE(DEVICE)
        )
    i_lut_985
        (
            .in_data({
                         in_data[723],
                         in_data[442],
                         in_data[2],
                         in_data[192],
                         in_data[255],
                         in_data[99]
                    }),
            .out_data(lut_985_out)
        );

reg   lut_985_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_985_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_985_ff <= lut_985_out;
    end
end

assign out_data[985] = lut_985_ff;




// LUT : 986

wire lut_986_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100011001111001000111101101011011111001101111001001011010100),
            .DEVICE(DEVICE)
        )
    i_lut_986
        (
            .in_data({
                         in_data[655],
                         in_data[123],
                         in_data[83],
                         in_data[690],
                         in_data[591],
                         in_data[726]
                    }),
            .out_data(lut_986_out)
        );

reg   lut_986_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_986_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_986_ff <= lut_986_out;
    end
end

assign out_data[986] = lut_986_ff;




// LUT : 987

wire lut_987_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010111001111101110000011101011000111000111110011001100011010),
            .DEVICE(DEVICE)
        )
    i_lut_987
        (
            .in_data({
                         in_data[353],
                         in_data[267],
                         in_data[364],
                         in_data[476],
                         in_data[209],
                         in_data[717]
                    }),
            .out_data(lut_987_out)
        );

reg   lut_987_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_987_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_987_ff <= lut_987_out;
    end
end

assign out_data[987] = lut_987_ff;




// LUT : 988

wire lut_988_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000100110100011110101001001011011011011001101111010001010010),
            .DEVICE(DEVICE)
        )
    i_lut_988
        (
            .in_data({
                         in_data[534],
                         in_data[393],
                         in_data[673],
                         in_data[681],
                         in_data[23],
                         in_data[51]
                    }),
            .out_data(lut_988_out)
        );

reg   lut_988_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_988_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_988_ff <= lut_988_out;
    end
end

assign out_data[988] = lut_988_ff;




// LUT : 989

wire lut_989_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010110011101100010000001111011100010110001001001001100010010001),
            .DEVICE(DEVICE)
        )
    i_lut_989
        (
            .in_data({
                         in_data[274],
                         in_data[74],
                         in_data[310],
                         in_data[615],
                         in_data[705],
                         in_data[410]
                    }),
            .out_data(lut_989_out)
        );

reg   lut_989_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_989_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_989_ff <= lut_989_out;
    end
end

assign out_data[989] = lut_989_ff;




// LUT : 990

wire lut_990_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011011110111110011111011111011101110100110111111010101011101010),
            .DEVICE(DEVICE)
        )
    i_lut_990
        (
            .in_data({
                         in_data[594],
                         in_data[36],
                         in_data[320],
                         in_data[294],
                         in_data[545],
                         in_data[251]
                    }),
            .out_data(lut_990_out)
        );

reg   lut_990_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_990_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_990_ff <= lut_990_out;
    end
end

assign out_data[990] = lut_990_ff;




// LUT : 991

wire lut_991_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010010000111101000111110111100000100110011101001010001011111),
            .DEVICE(DEVICE)
        )
    i_lut_991
        (
            .in_data({
                         in_data[109],
                         in_data[379],
                         in_data[417],
                         in_data[163],
                         in_data[713],
                         in_data[273]
                    }),
            .out_data(lut_991_out)
        );

reg   lut_991_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_991_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_991_ff <= lut_991_out;
    end
end

assign out_data[991] = lut_991_ff;




// LUT : 992

wire lut_992_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010011011010001000000000101000010110101110110001101001010001111),
            .DEVICE(DEVICE)
        )
    i_lut_992
        (
            .in_data({
                         in_data[256],
                         in_data[169],
                         in_data[321],
                         in_data[140],
                         in_data[355],
                         in_data[230]
                    }),
            .out_data(lut_992_out)
        );

reg   lut_992_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_992_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_992_ff <= lut_992_out;
    end
end

assign out_data[992] = lut_992_ff;




// LUT : 993

wire lut_993_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111010001000100001001010011101010011100100011100101010),
            .DEVICE(DEVICE)
        )
    i_lut_993
        (
            .in_data({
                         in_data[562],
                         in_data[701],
                         in_data[386],
                         in_data[727],
                         in_data[555],
                         in_data[730]
                    }),
            .out_data(lut_993_out)
        );

reg   lut_993_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_993_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_993_ff <= lut_993_out;
    end
end

assign out_data[993] = lut_993_ff;




// LUT : 994

wire lut_994_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100010111000101011100000100000000110111001000110011111100101010),
            .DEVICE(DEVICE)
        )
    i_lut_994
        (
            .in_data({
                         in_data[779],
                         in_data[190],
                         in_data[304],
                         in_data[116],
                         in_data[448],
                         in_data[610]
                    }),
            .out_data(lut_994_out)
        );

reg   lut_994_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_994_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_994_ff <= lut_994_out;
    end
end

assign out_data[994] = lut_994_ff;




// LUT : 995

wire lut_995_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100011101100101000111010100100011001000010011010100110010000000),
            .DEVICE(DEVICE)
        )
    i_lut_995
        (
            .in_data({
                         in_data[142],
                         in_data[481],
                         in_data[368],
                         in_data[463],
                         in_data[58],
                         in_data[497]
                    }),
            .out_data(lut_995_out)
        );

reg   lut_995_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_995_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_995_ff <= lut_995_out;
    end
end

assign out_data[995] = lut_995_ff;




// LUT : 996

wire lut_996_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111110000101101100011010111011000001100101001101110011010001),
            .DEVICE(DEVICE)
        )
    i_lut_996
        (
            .in_data({
                         in_data[675],
                         in_data[61],
                         in_data[453],
                         in_data[19],
                         in_data[643],
                         in_data[752]
                    }),
            .out_data(lut_996_out)
        );

reg   lut_996_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_996_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_996_ff <= lut_996_out;
    end
end

assign out_data[996] = lut_996_ff;




// LUT : 997

wire lut_997_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011000000000100100111010000010011110000000110010001001000001),
            .DEVICE(DEVICE)
        )
    i_lut_997
        (
            .in_data({
                         in_data[563],
                         in_data[272],
                         in_data[557],
                         in_data[301],
                         in_data[627],
                         in_data[735]
                    }),
            .out_data(lut_997_out)
        );

reg   lut_997_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_997_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_997_ff <= lut_997_out;
    end
end

assign out_data[997] = lut_997_ff;




// LUT : 998

wire lut_998_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110101110111010100010111001101010011110100100111110101111101),
            .DEVICE(DEVICE)
        )
    i_lut_998
        (
            .in_data({
                         in_data[220],
                         in_data[156],
                         in_data[344],
                         in_data[200],
                         in_data[186],
                         in_data[765]
                    }),
            .out_data(lut_998_out)
        );

reg   lut_998_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_998_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_998_ff <= lut_998_out;
    end
end

assign out_data[998] = lut_998_ff;




// LUT : 999

wire lut_999_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101011011011000011110100010010000101011011111111000001001010000),
            .DEVICE(DEVICE)
        )
    i_lut_999
        (
            .in_data({
                         in_data[559],
                         in_data[443],
                         in_data[227],
                         in_data[572],
                         in_data[548],
                         in_data[590]
                    }),
            .out_data(lut_999_out)
        );

reg   lut_999_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_999_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_999_ff <= lut_999_out;
    end
end

assign out_data[999] = lut_999_ff;




// LUT : 1000

wire lut_1000_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011010111110000101100011100000010101100111111111000000001110101),
            .DEVICE(DEVICE)
        )
    i_lut_1000
        (
            .in_data({
                         in_data[37],
                         in_data[523],
                         in_data[188],
                         in_data[518],
                         in_data[305],
                         in_data[580]
                    }),
            .out_data(lut_1000_out)
        );

reg   lut_1000_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1000_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1000_ff <= lut_1000_out;
    end
end

assign out_data[1000] = lut_1000_ff;




// LUT : 1001

wire lut_1001_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000111111111011010101111111101111111010100110111011100000011),
            .DEVICE(DEVICE)
        )
    i_lut_1001
        (
            .in_data({
                         in_data[749],
                         in_data[264],
                         in_data[474],
                         in_data[401],
                         in_data[324],
                         in_data[318]
                    }),
            .out_data(lut_1001_out)
        );

reg   lut_1001_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1001_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1001_ff <= lut_1001_out;
    end
end

assign out_data[1001] = lut_1001_ff;




// LUT : 1002

wire lut_1002_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100101011111000001100011001111000001100100110000010001110011),
            .DEVICE(DEVICE)
        )
    i_lut_1002
        (
            .in_data({
                         in_data[438],
                         in_data[671],
                         in_data[361],
                         in_data[495],
                         in_data[432],
                         in_data[266]
                    }),
            .out_data(lut_1002_out)
        );

reg   lut_1002_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1002_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1002_ff <= lut_1002_out;
    end
end

assign out_data[1002] = lut_1002_ff;




// LUT : 1003

wire lut_1003_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010111011101111101111111100001111101111111111101100110001010),
            .DEVICE(DEVICE)
        )
    i_lut_1003
        (
            .in_data({
                         in_data[648],
                         in_data[402],
                         in_data[662],
                         in_data[656],
                         in_data[325],
                         in_data[672]
                    }),
            .out_data(lut_1003_out)
        );

reg   lut_1003_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1003_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1003_ff <= lut_1003_out;
    end
end

assign out_data[1003] = lut_1003_ff;




// LUT : 1004

wire lut_1004_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000000010000000111010000111101001111001011101111111100101110),
            .DEVICE(DEVICE)
        )
    i_lut_1004
        (
            .in_data({
                         in_data[430],
                         in_data[338],
                         in_data[456],
                         in_data[659],
                         in_data[541],
                         in_data[136]
                    }),
            .out_data(lut_1004_out)
        );

reg   lut_1004_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1004_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1004_ff <= lut_1004_out;
    end
end

assign out_data[1004] = lut_1004_ff;




// LUT : 1005

wire lut_1005_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111101001111111110111111111110101011101010101010101111111111),
            .DEVICE(DEVICE)
        )
    i_lut_1005
        (
            .in_data({
                         in_data[144],
                         in_data[300],
                         in_data[285],
                         in_data[494],
                         in_data[356],
                         in_data[553]
                    }),
            .out_data(lut_1005_out)
        );

reg   lut_1005_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1005_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1005_ff <= lut_1005_out;
    end
end

assign out_data[1005] = lut_1005_ff;




// LUT : 1006

wire lut_1006_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110000001010111100001101010011110110010100110001011001100111100),
            .DEVICE(DEVICE)
        )
    i_lut_1006
        (
            .in_data({
                         in_data[778],
                         in_data[508],
                         in_data[704],
                         in_data[745],
                         in_data[12],
                         in_data[270]
                    }),
            .out_data(lut_1006_out)
        );

reg   lut_1006_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1006_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1006_ff <= lut_1006_out;
    end
end

assign out_data[1006] = lut_1006_ff;




// LUT : 1007

wire lut_1007_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001011111100100000100111000101010101001101010000111101101110111),
            .DEVICE(DEVICE)
        )
    i_lut_1007
        (
            .in_data({
                         in_data[689],
                         in_data[739],
                         in_data[677],
                         in_data[236],
                         in_data[15],
                         in_data[52]
                    }),
            .out_data(lut_1007_out)
        );

reg   lut_1007_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1007_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1007_ff <= lut_1007_out;
    end
end

assign out_data[1007] = lut_1007_ff;




// LUT : 1008

wire lut_1008_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001110010000101000101100111000010101011110100010100010001101),
            .DEVICE(DEVICE)
        )
    i_lut_1008
        (
            .in_data({
                         in_data[31],
                         in_data[641],
                         in_data[105],
                         in_data[247],
                         in_data[381],
                         in_data[782]
                    }),
            .out_data(lut_1008_out)
        );

reg   lut_1008_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1008_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1008_ff <= lut_1008_out;
    end
end

assign out_data[1008] = lut_1008_ff;




// LUT : 1009

wire lut_1009_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000001110111000011011011101111111000111100111000110000010001),
            .DEVICE(DEVICE)
        )
    i_lut_1009
        (
            .in_data({
                         in_data[245],
                         in_data[466],
                         in_data[632],
                         in_data[158],
                         in_data[168],
                         in_data[151]
                    }),
            .out_data(lut_1009_out)
        );

reg   lut_1009_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1009_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1009_ff <= lut_1009_out;
    end
end

assign out_data[1009] = lut_1009_ff;




// LUT : 1010

wire lut_1010_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101111111111100000010011111100001110110101011011001100110101),
            .DEVICE(DEVICE)
        )
    i_lut_1010
        (
            .in_data({
                         in_data[653],
                         in_data[759],
                         in_data[281],
                         in_data[288],
                         in_data[6],
                         in_data[85]
                    }),
            .out_data(lut_1010_out)
        );

reg   lut_1010_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1010_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1010_ff <= lut_1010_out;
    end
end

assign out_data[1010] = lut_1010_ff;




// LUT : 1011

wire lut_1011_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111101000001100000000010001000111010000110111111010010011101100),
            .DEVICE(DEVICE)
        )
    i_lut_1011
        (
            .in_data({
                         in_data[748],
                         in_data[183],
                         in_data[291],
                         in_data[10],
                         in_data[524],
                         in_data[384]
                    }),
            .out_data(lut_1011_out)
        );

reg   lut_1011_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1011_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1011_ff <= lut_1011_out;
    end
end

assign out_data[1011] = lut_1011_ff;




// LUT : 1012

wire lut_1012_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011100110011010010011011001111011010100000001110000101000101),
            .DEVICE(DEVICE)
        )
    i_lut_1012
        (
            .in_data({
                         in_data[57],
                         in_data[529],
                         in_data[124],
                         in_data[29],
                         in_data[510],
                         in_data[640]
                    }),
            .out_data(lut_1012_out)
        );

reg   lut_1012_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1012_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1012_ff <= lut_1012_out;
    end
end

assign out_data[1012] = lut_1012_ff;




// LUT : 1013

wire lut_1013_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001110101111010011011101110010001111100101111110111111111100),
            .DEVICE(DEVICE)
        )
    i_lut_1013
        (
            .in_data({
                         in_data[493],
                         in_data[108],
                         in_data[606],
                         in_data[279],
                         in_data[303],
                         in_data[351]
                    }),
            .out_data(lut_1013_out)
        );

reg   lut_1013_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1013_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1013_ff <= lut_1013_out;
    end
end

assign out_data[1013] = lut_1013_ff;




// LUT : 1014

wire lut_1014_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100011111001001101111100100001001000001100110010001011110010),
            .DEVICE(DEVICE)
        )
    i_lut_1014
        (
            .in_data({
                         in_data[362],
                         in_data[736],
                         in_data[638],
                         in_data[290],
                         in_data[688],
                         in_data[265]
                    }),
            .out_data(lut_1014_out)
        );

reg   lut_1014_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1014_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1014_ff <= lut_1014_out;
    end
end

assign out_data[1014] = lut_1014_ff;




// LUT : 1015

wire lut_1015_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000000100111010110101101110110101101011010110111111111011101),
            .DEVICE(DEVICE)
        )
    i_lut_1015
        (
            .in_data({
                         in_data[629],
                         in_data[605],
                         in_data[342],
                         in_data[289],
                         in_data[354],
                         in_data[13]
                    }),
            .out_data(lut_1015_out)
        );

reg   lut_1015_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1015_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1015_ff <= lut_1015_out;
    end
end

assign out_data[1015] = lut_1015_ff;




// LUT : 1016

wire lut_1016_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001000000100101010000001000010011010010101001011111001000100101),
            .DEVICE(DEVICE)
        )
    i_lut_1016
        (
            .in_data({
                         in_data[185],
                         in_data[436],
                         in_data[623],
                         in_data[366],
                         in_data[491],
                         in_data[418]
                    }),
            .out_data(lut_1016_out)
        );

reg   lut_1016_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1016_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1016_ff <= lut_1016_out;
    end
end

assign out_data[1016] = lut_1016_ff;




// LUT : 1017

wire lut_1017_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110000100100001001011010010101111111011010000010011100101000001),
            .DEVICE(DEVICE)
        )
    i_lut_1017
        (
            .in_data({
                         in_data[692],
                         in_data[539],
                         in_data[101],
                         in_data[240],
                         in_data[746],
                         in_data[308]
                    }),
            .out_data(lut_1017_out)
        );

reg   lut_1017_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1017_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1017_ff <= lut_1017_out;
    end
end

assign out_data[1017] = lut_1017_ff;




// LUT : 1018

wire lut_1018_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110010000000111011010111000000111100010010000000110010001100),
            .DEVICE(DEVICE)
        )
    i_lut_1018
        (
            .in_data({
                         in_data[250],
                         in_data[126],
                         in_data[441],
                         in_data[8],
                         in_data[568],
                         in_data[154]
                    }),
            .out_data(lut_1018_out)
        );

reg   lut_1018_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1018_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1018_ff <= lut_1018_out;
    end
end

assign out_data[1018] = lut_1018_ff;




// LUT : 1019

wire lut_1019_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011001011111011000010101110101000010011100110110101101100101),
            .DEVICE(DEVICE)
        )
    i_lut_1019
        (
            .in_data({
                         in_data[551],
                         in_data[44],
                         in_data[1],
                         in_data[98],
                         in_data[218],
                         in_data[298]
                    }),
            .out_data(lut_1019_out)
        );

reg   lut_1019_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1019_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1019_ff <= lut_1019_out;
    end
end

assign out_data[1019] = lut_1019_ff;




// LUT : 1020

wire lut_1020_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011100100100010100010101011110100000111101101010001100000110),
            .DEVICE(DEVICE)
        )
    i_lut_1020
        (
            .in_data({
                         in_data[161],
                         in_data[770],
                         in_data[392],
                         in_data[24],
                         in_data[306],
                         in_data[191]
                    }),
            .out_data(lut_1020_out)
        );

reg   lut_1020_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1020_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1020_ff <= lut_1020_out;
    end
end

assign out_data[1020] = lut_1020_ff;




// LUT : 1021

wire lut_1021_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010100000001111000000001000111001001000001011100000000001000110),
            .DEVICE(DEVICE)
        )
    i_lut_1021
        (
            .in_data({
                         in_data[737],
                         in_data[760],
                         in_data[498],
                         in_data[248],
                         in_data[374],
                         in_data[549]
                    }),
            .out_data(lut_1021_out)
        );

reg   lut_1021_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1021_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1021_ff <= lut_1021_out;
    end
end

assign out_data[1021] = lut_1021_ff;




// LUT : 1022

wire lut_1022_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110001110100011110010111111101100011100011001001011101011111),
            .DEVICE(DEVICE)
        )
    i_lut_1022
        (
            .in_data({
                         in_data[94],
                         in_data[634],
                         in_data[695],
                         in_data[276],
                         in_data[519],
                         in_data[42]
                    }),
            .out_data(lut_1022_out)
        );

reg   lut_1022_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1022_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1022_ff <= lut_1022_out;
    end
end

assign out_data[1022] = lut_1022_ff;




// LUT : 1023

wire lut_1023_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101010110111110110101000110110100001100001010000110110000101),
            .DEVICE(DEVICE)
        )
    i_lut_1023
        (
            .in_data({
                         in_data[334],
                         in_data[257],
                         in_data[397],
                         in_data[358],
                         in_data[462],
                         in_data[774]
                    }),
            .out_data(lut_1023_out)
        );

reg   lut_1023_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1023_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1023_ff <= lut_1023_out;
    end
end

assign out_data[1023] = lut_1023_ff;



endmodule



module MnistStochasticLut6Mlp_sub1
        #(
            parameter DEVICE = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [1023:0]  in_data,
            output wire [359:0]  out_data
        );


// LUT : 0

wire lut_0_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110111111011111110011011111111111101111100001010100110111),
            .DEVICE(DEVICE)
        )
    i_lut_0
        (
            .in_data({
                         in_data[111],
                         in_data[736],
                         in_data[420],
                         in_data[803],
                         in_data[302],
                         in_data[531]
                    }),
            .out_data(lut_0_out)
        );

reg   lut_0_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_0_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_0_ff <= lut_0_out;
    end
end

assign out_data[0] = lut_0_ff;




// LUT : 1

wire lut_1_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000001000000010000000100000001100111011100000111011001110),
            .DEVICE(DEVICE)
        )
    i_lut_1
        (
            .in_data({
                         in_data[20],
                         in_data[400],
                         in_data[203],
                         in_data[529],
                         in_data[832],
                         in_data[812]
                    }),
            .out_data(lut_1_out)
        );

reg   lut_1_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1_ff <= lut_1_out;
    end
end

assign out_data[1] = lut_1_ff;




// LUT : 2

wire lut_2_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111110011011111111110011001101111101001010100),
            .DEVICE(DEVICE)
        )
    i_lut_2
        (
            .in_data({
                         in_data[898],
                         in_data[148],
                         in_data[725],
                         in_data[692],
                         in_data[677],
                         in_data[620]
                    }),
            .out_data(lut_2_out)
        );

reg   lut_2_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_2_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_2_ff <= lut_2_out;
    end
end

assign out_data[2] = lut_2_ff;




// LUT : 3

wire lut_3_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111101111111101111001111111010001110011110001101111001111),
            .DEVICE(DEVICE)
        )
    i_lut_3
        (
            .in_data({
                         in_data[330],
                         in_data[606],
                         in_data[98],
                         in_data[501],
                         in_data[44],
                         in_data[663]
                    }),
            .out_data(lut_3_out)
        );

reg   lut_3_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_3_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_3_ff <= lut_3_out;
    end
end

assign out_data[3] = lut_3_ff;




// LUT : 4

wire lut_4_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111011111110001111111111111111011111111111100110111),
            .DEVICE(DEVICE)
        )
    i_lut_4
        (
            .in_data({
                         in_data[932],
                         in_data[967],
                         in_data[939],
                         in_data[129],
                         in_data[742],
                         in_data[334]
                    }),
            .out_data(lut_4_out)
        );

reg   lut_4_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_4_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_4_ff <= lut_4_out;
    end
end

assign out_data[4] = lut_4_ff;




// LUT : 5

wire lut_5_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111111111111111011111111100111000101010100001100110001011001),
            .DEVICE(DEVICE)
        )
    i_lut_5
        (
            .in_data({
                         in_data[574],
                         in_data[419],
                         in_data[699],
                         in_data[193],
                         in_data[298],
                         in_data[771]
                    }),
            .out_data(lut_5_out)
        );

reg   lut_5_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_5_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_5_ff <= lut_5_out;
    end
end

assign out_data[5] = lut_5_ff;




// LUT : 6

wire lut_6_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010011111100000000000000000011111101111010001100110110000101),
            .DEVICE(DEVICE)
        )
    i_lut_6
        (
            .in_data({
                         in_data[966],
                         in_data[359],
                         in_data[580],
                         in_data[999],
                         in_data[608],
                         in_data[783]
                    }),
            .out_data(lut_6_out)
        );

reg   lut_6_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_6_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_6_ff <= lut_6_out;
    end
end

assign out_data[6] = lut_6_ff;




// LUT : 7

wire lut_7_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001000000010100100000001001000000000000000101001000000100),
            .DEVICE(DEVICE)
        )
    i_lut_7
        (
            .in_data({
                         in_data[338],
                         in_data[936],
                         in_data[424],
                         in_data[502],
                         in_data[320],
                         in_data[696]
                    }),
            .out_data(lut_7_out)
        );

reg   lut_7_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_7_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_7_ff <= lut_7_out;
    end
end

assign out_data[7] = lut_7_ff;




// LUT : 8

wire lut_8_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111110110111011111111011101110111111100010111111110000110011),
            .DEVICE(DEVICE)
        )
    i_lut_8
        (
            .in_data({
                         in_data[394],
                         in_data[101],
                         in_data[512],
                         in_data[490],
                         in_data[480],
                         in_data[433]
                    }),
            .out_data(lut_8_out)
        );

reg   lut_8_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_8_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_8_ff <= lut_8_out;
    end
end

assign out_data[8] = lut_8_ff;




// LUT : 9

wire lut_9_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001101101101111111111101111111100010000000000111111001000101011),
            .DEVICE(DEVICE)
        )
    i_lut_9
        (
            .in_data({
                         in_data[882],
                         in_data[322],
                         in_data[745],
                         in_data[472],
                         in_data[141],
                         in_data[972]
                    }),
            .out_data(lut_9_out)
        );

reg   lut_9_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_9_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_9_ff <= lut_9_out;
    end
end

assign out_data[9] = lut_9_ff;




// LUT : 10

wire lut_10_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001000000000000000010000110000000011000011000000011100001111),
            .DEVICE(DEVICE)
        )
    i_lut_10
        (
            .in_data({
                         in_data[561],
                         in_data[629],
                         in_data[252],
                         in_data[522],
                         in_data[983],
                         in_data[296]
                    }),
            .out_data(lut_10_out)
        );

reg   lut_10_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_10_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_10_ff <= lut_10_out;
    end
end

assign out_data[10] = lut_10_ff;




// LUT : 11

wire lut_11_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010011011101110100001011100000111000110111101101001111110111111),
            .DEVICE(DEVICE)
        )
    i_lut_11
        (
            .in_data({
                         in_data[125],
                         in_data[820],
                         in_data[850],
                         in_data[560],
                         in_data[53],
                         in_data[689]
                    }),
            .out_data(lut_11_out)
        );

reg   lut_11_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_11_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_11_ff <= lut_11_out;
    end
end

assign out_data[11] = lut_11_ff;




// LUT : 12

wire lut_12_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010111100101111000111110111101100001011000011110000110100111101),
            .DEVICE(DEVICE)
        )
    i_lut_12
        (
            .in_data({
                         in_data[123],
                         in_data[147],
                         in_data[340],
                         in_data[602],
                         in_data[171],
                         in_data[789]
                    }),
            .out_data(lut_12_out)
        );

reg   lut_12_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_12_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_12_ff <= lut_12_out;
    end
end

assign out_data[12] = lut_12_ff;




// LUT : 13

wire lut_13_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110010000011000011111101111100000101101100000000111100000111),
            .DEVICE(DEVICE)
        )
    i_lut_13
        (
            .in_data({
                         in_data[513],
                         in_data[990],
                         in_data[840],
                         in_data[168],
                         in_data[128],
                         in_data[232]
                    }),
            .out_data(lut_13_out)
        );

reg   lut_13_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_13_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_13_ff <= lut_13_out;
    end
end

assign out_data[13] = lut_13_ff;




// LUT : 14

wire lut_14_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001011010111111101100001110011001010100101111101011001011110010),
            .DEVICE(DEVICE)
        )
    i_lut_14
        (
            .in_data({
                         in_data[526],
                         in_data[276],
                         in_data[352],
                         in_data[844],
                         in_data[993],
                         in_data[970]
                    }),
            .out_data(lut_14_out)
        );

reg   lut_14_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_14_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_14_ff <= lut_14_out;
    end
end

assign out_data[14] = lut_14_ff;




// LUT : 15

wire lut_15_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111000000001110101011111111111111111110000011111110),
            .DEVICE(DEVICE)
        )
    i_lut_15
        (
            .in_data({
                         in_data[600],
                         in_data[79],
                         in_data[267],
                         in_data[804],
                         in_data[935],
                         in_data[701]
                    }),
            .out_data(lut_15_out)
        );

reg   lut_15_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_15_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_15_ff <= lut_15_out;
    end
end

assign out_data[15] = lut_15_ff;




// LUT : 16

wire lut_16_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000010011100101100000100110000011000000011110000000001001110),
            .DEVICE(DEVICE)
        )
    i_lut_16
        (
            .in_data({
                         in_data[353],
                         in_data[116],
                         in_data[337],
                         in_data[58],
                         in_data[97],
                         in_data[368]
                    }),
            .out_data(lut_16_out)
        );

reg   lut_16_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_16_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_16_ff <= lut_16_out;
    end
end

assign out_data[16] = lut_16_ff;




// LUT : 17

wire lut_17_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000010000000110100000101001000000100000001000101000011010000),
            .DEVICE(DEVICE)
        )
    i_lut_17
        (
            .in_data({
                         in_data[304],
                         in_data[221],
                         in_data[738],
                         in_data[481],
                         in_data[749],
                         in_data[77]
                    }),
            .out_data(lut_17_out)
        );

reg   lut_17_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_17_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_17_ff <= lut_17_out;
    end
end

assign out_data[17] = lut_17_ff;




// LUT : 18

wire lut_18_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111111111111100000111111111111011111111110111101111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_18
        (
            .in_data({
                         in_data[152],
                         in_data[805],
                         in_data[33],
                         in_data[946],
                         in_data[374],
                         in_data[506]
                    }),
            .out_data(lut_18_out)
        );

reg   lut_18_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_18_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_18_ff <= lut_18_out;
    end
end

assign out_data[18] = lut_18_ff;




// LUT : 19

wire lut_19_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101111100010111011001110111101010100111101001100110011001101),
            .DEVICE(DEVICE)
        )
    i_lut_19
        (
            .in_data({
                         in_data[605],
                         in_data[389],
                         in_data[565],
                         in_data[728],
                         in_data[365],
                         in_data[166]
                    }),
            .out_data(lut_19_out)
        );

reg   lut_19_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_19_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_19_ff <= lut_19_out;
    end
end

assign out_data[19] = lut_19_ff;




// LUT : 20

wire lut_20_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111111101100011001111100110011111111111111111111111110111101),
            .DEVICE(DEVICE)
        )
    i_lut_20
        (
            .in_data({
                         in_data[64],
                         in_data[852],
                         in_data[436],
                         in_data[427],
                         in_data[172],
                         in_data[393]
                    }),
            .out_data(lut_20_out)
        );

reg   lut_20_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_20_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_20_ff <= lut_20_out;
    end
end

assign out_data[20] = lut_20_ff;




// LUT : 21

wire lut_21_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000111111111111110110000000001000000110110000000001100000100),
            .DEVICE(DEVICE)
        )
    i_lut_21
        (
            .in_data({
                         in_data[54],
                         in_data[435],
                         in_data[549],
                         in_data[662],
                         in_data[928],
                         in_data[208]
                    }),
            .out_data(lut_21_out)
        );

reg   lut_21_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_21_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_21_ff <= lut_21_out;
    end
end

assign out_data[21] = lut_21_ff;




// LUT : 22

wire lut_22_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101111111110011110101101110111110011111111111101000111011101),
            .DEVICE(DEVICE)
        )
    i_lut_22
        (
            .in_data({
                         in_data[43],
                         in_data[107],
                         in_data[444],
                         in_data[628],
                         in_data[332],
                         in_data[431]
                    }),
            .out_data(lut_22_out)
        );

reg   lut_22_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_22_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_22_ff <= lut_22_out;
    end
end

assign out_data[22] = lut_22_ff;




// LUT : 23

wire lut_23_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001100101111000100011011111100110011001011110011001111111111),
            .DEVICE(DEVICE)
        )
    i_lut_23
        (
            .in_data({
                         in_data[648],
                         in_data[890],
                         in_data[924],
                         in_data[622],
                         in_data[788],
                         in_data[874]
                    }),
            .out_data(lut_23_out)
        );

reg   lut_23_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_23_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_23_ff <= lut_23_out;
    end
end

assign out_data[23] = lut_23_ff;




// LUT : 24

wire lut_24_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101011011111111111101111111111111010111111101111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_24
        (
            .in_data({
                         in_data[511],
                         in_data[155],
                         in_data[510],
                         in_data[724],
                         in_data[907],
                         in_data[269]
                    }),
            .out_data(lut_24_out)
        );

reg   lut_24_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_24_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_24_ff <= lut_24_out;
    end
end

assign out_data[24] = lut_24_ff;




// LUT : 25

wire lut_25_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010001000110000000000000011011000100100001001100000001000000),
            .DEVICE(DEVICE)
        )
    i_lut_25
        (
            .in_data({
                         in_data[63],
                         in_data[459],
                         in_data[504],
                         in_data[142],
                         in_data[923],
                         in_data[601]
                    }),
            .out_data(lut_25_out)
        );

reg   lut_25_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_25_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_25_ff <= lut_25_out;
    end
end

assign out_data[25] = lut_25_ff;




// LUT : 26

wire lut_26_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010011000010010101010001001101110110011111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_26
        (
            .in_data({
                         in_data[361],
                         in_data[236],
                         in_data[1013],
                         in_data[817],
                         in_data[179],
                         in_data[131]
                    }),
            .out_data(lut_26_out)
        );

reg   lut_26_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_26_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_26_ff <= lut_26_out;
    end
end

assign out_data[26] = lut_26_ff;




// LUT : 27

wire lut_27_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000011000111000001111100000000001000110011000100110011),
            .DEVICE(DEVICE)
        )
    i_lut_27
        (
            .in_data({
                         in_data[717],
                         in_data[793],
                         in_data[494],
                         in_data[223],
                         in_data[521],
                         in_data[432]
                    }),
            .out_data(lut_27_out)
        );

reg   lut_27_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_27_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_27_ff <= lut_27_out;
    end
end

assign out_data[27] = lut_27_ff;




// LUT : 28

wire lut_28_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000011100000000000001010100000010100010001000100000100000101),
            .DEVICE(DEVICE)
        )
    i_lut_28
        (
            .in_data({
                         in_data[678],
                         in_data[774],
                         in_data[84],
                         in_data[634],
                         in_data[2],
                         in_data[528]
                    }),
            .out_data(lut_28_out)
        );

reg   lut_28_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_28_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_28_ff <= lut_28_out;
    end
end

assign out_data[28] = lut_28_ff;




// LUT : 29

wire lut_29_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001001111111000000000111101011111111111111111111001011110010),
            .DEVICE(DEVICE)
        )
    i_lut_29
        (
            .in_data({
                         in_data[706],
                         in_data[130],
                         in_data[959],
                         in_data[488],
                         in_data[786],
                         in_data[870]
                    }),
            .out_data(lut_29_out)
        );

reg   lut_29_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_29_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_29_ff <= lut_29_out;
    end
end

assign out_data[29] = lut_29_ff;




// LUT : 30

wire lut_30_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001010000100001010101000010001101101001011100100011001011100110),
            .DEVICE(DEVICE)
        )
    i_lut_30
        (
            .in_data({
                         in_data[286],
                         in_data[920],
                         in_data[415],
                         in_data[333],
                         in_data[151],
                         in_data[576]
                    }),
            .out_data(lut_30_out)
        );

reg   lut_30_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_30_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_30_ff <= lut_30_out;
    end
end

assign out_data[30] = lut_30_ff;




// LUT : 31

wire lut_31_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111110001100111111111100111111011111110011000000011111001111),
            .DEVICE(DEVICE)
        )
    i_lut_31
        (
            .in_data({
                         in_data[228],
                         in_data[408],
                         in_data[160],
                         in_data[437],
                         in_data[779],
                         in_data[649]
                    }),
            .out_data(lut_31_out)
        );

reg   lut_31_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_31_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_31_ff <= lut_31_out;
    end
end

assign out_data[31] = lut_31_ff;




// LUT : 32

wire lut_32_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111100000010111011111110111110000001000001111110111111010),
            .DEVICE(DEVICE)
        )
    i_lut_32
        (
            .in_data({
                         in_data[60],
                         in_data[465],
                         in_data[294],
                         in_data[402],
                         in_data[229],
                         in_data[914]
                    }),
            .out_data(lut_32_out)
        );

reg   lut_32_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_32_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_32_ff <= lut_32_out;
    end
end

assign out_data[32] = lut_32_ff;




// LUT : 33

wire lut_33_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001001100000001110100000000000010000000000100011001100000000),
            .DEVICE(DEVICE)
        )
    i_lut_33
        (
            .in_data({
                         in_data[787],
                         in_data[943],
                         in_data[318],
                         in_data[958],
                         in_data[912],
                         in_data[39]
                    }),
            .out_data(lut_33_out)
        );

reg   lut_33_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_33_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_33_ff <= lut_33_out;
    end
end

assign out_data[33] = lut_33_ff;




// LUT : 34

wire lut_34_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001010111111101010100010101110111000110111001101101011010010),
            .DEVICE(DEVICE)
        )
    i_lut_34
        (
            .in_data({
                         in_data[806],
                         in_data[809],
                         in_data[76],
                         in_data[863],
                         in_data[756],
                         in_data[113]
                    }),
            .out_data(lut_34_out)
        );

reg   lut_34_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_34_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_34_ff <= lut_34_out;
    end
end

assign out_data[34] = lut_34_ff;




// LUT : 35

wire lut_35_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101111110011111100111111111110110010011101100111001000110110),
            .DEVICE(DEVICE)
        )
    i_lut_35
        (
            .in_data({
                         in_data[190],
                         in_data[934],
                         in_data[209],
                         in_data[418],
                         in_data[92],
                         in_data[590]
                    }),
            .out_data(lut_35_out)
        );

reg   lut_35_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_35_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_35_ff <= lut_35_out;
    end
end

assign out_data[35] = lut_35_ff;




// LUT : 36

wire lut_36_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111110111010101011111111100110000001100000011001111110011),
            .DEVICE(DEVICE)
        )
    i_lut_36
        (
            .in_data({
                         in_data[642],
                         in_data[652],
                         in_data[370],
                         in_data[367],
                         in_data[571],
                         in_data[796]
                    }),
            .out_data(lut_36_out)
        );

reg   lut_36_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_36_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_36_ff <= lut_36_out;
    end
end

assign out_data[36] = lut_36_ff;




// LUT : 37

wire lut_37_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001000101011001000110011101111100000010000100011010001000000),
            .DEVICE(DEVICE)
        )
    i_lut_37
        (
            .in_data({
                         in_data[22],
                         in_data[611],
                         in_data[482],
                         in_data[399],
                         in_data[478],
                         in_data[134]
                    }),
            .out_data(lut_37_out)
        );

reg   lut_37_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_37_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_37_ff <= lut_37_out;
    end
end

assign out_data[37] = lut_37_ff;




// LUT : 38

wire lut_38_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000010101011000000000000000000000001001100110011000001000000),
            .DEVICE(DEVICE)
        )
    i_lut_38
        (
            .in_data({
                         in_data[818],
                         in_data[851],
                         in_data[886],
                         in_data[491],
                         in_data[570],
                         in_data[487]
                    }),
            .out_data(lut_38_out)
        );

reg   lut_38_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_38_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_38_ff <= lut_38_out;
    end
end

assign out_data[38] = lut_38_ff;




// LUT : 39

wire lut_39_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111011111010000111110111101010100010101000000000001000100),
            .DEVICE(DEVICE)
        )
    i_lut_39
        (
            .in_data({
                         in_data[666],
                         in_data[916],
                         in_data[114],
                         in_data[894],
                         in_data[336],
                         in_data[328]
                    }),
            .out_data(lut_39_out)
        );

reg   lut_39_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_39_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_39_ff <= lut_39_out;
    end
end

assign out_data[39] = lut_39_ff;




// LUT : 40

wire lut_40_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111101100011111111110110011111111111111100110111100000000),
            .DEVICE(DEVICE)
        )
    i_lut_40
        (
            .in_data({
                         in_data[364],
                         in_data[173],
                         in_data[326],
                         in_data[603],
                         in_data[1021],
                         in_data[982]
                    }),
            .out_data(lut_40_out)
        );

reg   lut_40_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_40_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_40_ff <= lut_40_out;
    end
end

assign out_data[40] = lut_40_ff;




// LUT : 41

wire lut_41_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111111001110110111111110101011111111111110111111111111111010),
            .DEVICE(DEVICE)
        )
    i_lut_41
        (
            .in_data({
                         in_data[210],
                         in_data[452],
                         in_data[473],
                         in_data[913],
                         in_data[956],
                         in_data[174]
                    }),
            .out_data(lut_41_out)
        );

reg   lut_41_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_41_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_41_ff <= lut_41_out;
    end
end

assign out_data[41] = lut_41_ff;




// LUT : 42

wire lut_42_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110010000000111111111111101011111111111111101111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_42
        (
            .in_data({
                         in_data[238],
                         in_data[548],
                         in_data[887],
                         in_data[858],
                         in_data[635],
                         in_data[811]
                    }),
            .out_data(lut_42_out)
        );

reg   lut_42_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_42_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_42_ff <= lut_42_out;
    end
end

assign out_data[42] = lut_42_ff;




// LUT : 43

wire lut_43_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111110111111010111110011111110111010101110111011111110111011),
            .DEVICE(DEVICE)
        )
    i_lut_43
        (
            .in_data({
                         in_data[271],
                         in_data[138],
                         in_data[987],
                         in_data[307],
                         in_data[964],
                         in_data[976]
                    }),
            .out_data(lut_43_out)
        );

reg   lut_43_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_43_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_43_ff <= lut_43_out;
    end
end

assign out_data[43] = lut_43_ff;




// LUT : 44

wire lut_44_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000000000000000001100000000011001100000000001000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_44
        (
            .in_data({
                         in_data[578],
                         in_data[896],
                         in_data[937],
                         in_data[640],
                         in_data[95],
                         in_data[873]
                    }),
            .out_data(lut_44_out)
        );

reg   lut_44_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_44_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_44_ff <= lut_44_out;
    end
end

assign out_data[44] = lut_44_ff;




// LUT : 45

wire lut_45_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111100001111100111111111111111111111110011110100),
            .DEVICE(DEVICE)
        )
    i_lut_45
        (
            .in_data({
                         in_data[373],
                         in_data[973],
                         in_data[1009],
                         in_data[671],
                         in_data[299],
                         in_data[460]
                    }),
            .out_data(lut_45_out)
        );

reg   lut_45_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_45_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_45_ff <= lut_45_out;
    end
end

assign out_data[45] = lut_45_ff;




// LUT : 46

wire lut_46_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100101111001111110010101110101000000010010011111100001011110010),
            .DEVICE(DEVICE)
        )
    i_lut_46
        (
            .in_data({
                         in_data[509],
                         in_data[170],
                         in_data[750],
                         in_data[905],
                         in_data[888],
                         in_data[540]
                    }),
            .out_data(lut_46_out)
        );

reg   lut_46_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_46_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_46_ff <= lut_46_out;
    end
end

assign out_data[46] = lut_46_ff;




// LUT : 47

wire lut_47_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000100011111001101110000111111111101011101010001000100000010),
            .DEVICE(DEVICE)
        )
    i_lut_47
        (
            .in_data({
                         in_data[297],
                         in_data[70],
                         in_data[633],
                         in_data[288],
                         in_data[849],
                         in_data[83]
                    }),
            .out_data(lut_47_out)
        );

reg   lut_47_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_47_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_47_ff <= lut_47_out;
    end
end

assign out_data[47] = lut_47_ff;




// LUT : 48

wire lut_48_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001000100000001000000000000000100010101000000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_48
        (
            .in_data({
                         in_data[930],
                         in_data[184],
                         in_data[117],
                         in_data[303],
                         in_data[827],
                         in_data[651]
                    }),
            .out_data(lut_48_out)
        );

reg   lut_48_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_48_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_48_ff <= lut_48_out;
    end
end

assign out_data[48] = lut_48_ff;




// LUT : 49

wire lut_49_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000101000000010000011000000000000001111000011110000),
            .DEVICE(DEVICE)
        )
    i_lut_49
        (
            .in_data({
                         in_data[950],
                         in_data[375],
                         in_data[163],
                         in_data[856],
                         in_data[822],
                         in_data[56]
                    }),
            .out_data(lut_49_out)
        );

reg   lut_49_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_49_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_49_ff <= lut_49_out;
    end
end

assign out_data[49] = lut_49_ff;




// LUT : 50

wire lut_50_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110011001111111111101101111011101101110000101111011001011100),
            .DEVICE(DEVICE)
        )
    i_lut_50
        (
            .in_data({
                         in_data[306],
                         in_data[604],
                         in_data[277],
                         in_data[268],
                         in_data[458],
                         in_data[627]
                    }),
            .out_data(lut_50_out)
        );

reg   lut_50_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_50_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_50_ff <= lut_50_out;
    end
end

assign out_data[50] = lut_50_ff;




// LUT : 51

wire lut_51_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101010100111101100000001000011111111111111111011011101101011),
            .DEVICE(DEVICE)
        )
    i_lut_51
        (
            .in_data({
                         in_data[589],
                         in_data[213],
                         in_data[797],
                         in_data[925],
                         in_data[566],
                         in_data[902]
                    }),
            .out_data(lut_51_out)
        );

reg   lut_51_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_51_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_51_ff <= lut_51_out;
    end
end

assign out_data[51] = lut_51_ff;




// LUT : 52

wire lut_52_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101001110000101010100010001100111010010100011110111011101111),
            .DEVICE(DEVICE)
        )
    i_lut_52
        (
            .in_data({
                         in_data[165],
                         in_data[572],
                         in_data[126],
                         in_data[638],
                         in_data[31],
                         in_data[423]
                    }),
            .out_data(lut_52_out)
        );

reg   lut_52_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_52_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_52_ff <= lut_52_out;
    end
end

assign out_data[52] = lut_52_ff;




// LUT : 53

wire lut_53_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111101101110111001111110111011011111111110111011111111101111101),
            .DEVICE(DEVICE)
        )
    i_lut_53
        (
            .in_data({
                         in_data[7],
                         in_data[667],
                         in_data[300],
                         in_data[564],
                         in_data[466],
                         in_data[895]
                    }),
            .out_data(lut_53_out)
        );

reg   lut_53_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_53_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_53_ff <= lut_53_out;
    end
end

assign out_data[53] = lut_53_ff;




// LUT : 54

wire lut_54_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001101100011111110011000101110110110110011111001101110010101001),
            .DEVICE(DEVICE)
        )
    i_lut_54
        (
            .in_data({
                         in_data[879],
                         in_data[313],
                         in_data[1020],
                         in_data[6],
                         in_data[537],
                         in_data[29]
                    }),
            .out_data(lut_54_out)
        );

reg   lut_54_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_54_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_54_ff <= lut_54_out;
    end
end

assign out_data[54] = lut_54_ff;




// LUT : 55

wire lut_55_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010000000101000001000000010000000100000011010000010000001100),
            .DEVICE(DEVICE)
        )
    i_lut_55
        (
            .in_data({
                         in_data[255],
                         in_data[938],
                         in_data[637],
                         in_data[527],
                         in_data[18],
                         in_data[467]
                    }),
            .out_data(lut_55_out)
        );

reg   lut_55_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_55_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_55_ff <= lut_55_out;
    end
end

assign out_data[55] = lut_55_ff;




// LUT : 56

wire lut_56_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111100101111111111110111101111111111001011111111111100111110),
            .DEVICE(DEVICE)
        )
    i_lut_56
        (
            .in_data({
                         in_data[729],
                         in_data[217],
                         in_data[106],
                         in_data[461],
                         in_data[759],
                         in_data[757]
                    }),
            .out_data(lut_56_out)
        );

reg   lut_56_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_56_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_56_ff <= lut_56_out;
    end
end

assign out_data[56] = lut_56_ff;




// LUT : 57

wire lut_57_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101011100000111110001101101101001011110110110101101001011011),
            .DEVICE(DEVICE)
        )
    i_lut_57
        (
            .in_data({
                         in_data[726],
                         in_data[146],
                         in_data[883],
                         in_data[242],
                         in_data[617],
                         in_data[650]
                    }),
            .out_data(lut_57_out)
        );

reg   lut_57_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_57_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_57_ff <= lut_57_out;
    end
end

assign out_data[57] = lut_57_ff;




// LUT : 58

wire lut_58_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111100000010011100001000000000000000000010000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_58
        (
            .in_data({
                         in_data[395],
                         in_data[158],
                         in_data[350],
                         in_data[957],
                         in_data[463],
                         in_data[778]
                    }),
            .out_data(lut_58_out)
        );

reg   lut_58_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_58_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_58_ff <= lut_58_out;
    end
end

assign out_data[58] = lut_58_ff;




// LUT : 59

wire lut_59_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000000011111000101010000011100010001000111010011011100001111),
            .DEVICE(DEVICE)
        )
    i_lut_59
        (
            .in_data({
                         in_data[655],
                         in_data[704],
                         in_data[746],
                         in_data[953],
                         in_data[777],
                         in_data[372]
                    }),
            .out_data(lut_59_out)
        );

reg   lut_59_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_59_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_59_ff <= lut_59_out;
    end
end

assign out_data[59] = lut_59_ff;




// LUT : 60

wire lut_60_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110111111101000011001101110011011101111111110001001010111011),
            .DEVICE(DEVICE)
        )
    i_lut_60
        (
            .in_data({
                         in_data[785],
                         in_data[703],
                         in_data[933],
                         in_data[665],
                         in_data[995],
                         in_data[291]
                    }),
            .out_data(lut_60_out)
        );

reg   lut_60_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_60_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_60_ff <= lut_60_out;
    end
end

assign out_data[60] = lut_60_ff;




// LUT : 61

wire lut_61_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001010001000001110101010100000000000000010000010100000101),
            .DEVICE(DEVICE)
        )
    i_lut_61
        (
            .in_data({
                         in_data[836],
                         in_data[290],
                         in_data[96],
                         in_data[247],
                         in_data[136],
                         in_data[544]
                    }),
            .out_data(lut_61_out)
        );

reg   lut_61_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_61_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_61_ff <= lut_61_out;
    end
end

assign out_data[61] = lut_61_ff;




// LUT : 62

wire lut_62_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000010110010100000001111001111100100011001100110000000100000101),
            .DEVICE(DEVICE)
        )
    i_lut_62
        (
            .in_data({
                         in_data[963],
                         in_data[497],
                         in_data[539],
                         in_data[360],
                         in_data[899],
                         in_data[455]
                    }),
            .out_data(lut_62_out)
        );

reg   lut_62_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_62_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_62_ff <= lut_62_out;
    end
end

assign out_data[62] = lut_62_ff;




// LUT : 63

wire lut_63_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000000000010010000000000000000000110100001111),
            .DEVICE(DEVICE)
        )
    i_lut_63
        (
            .in_data({
                         in_data[609],
                         in_data[686],
                         in_data[102],
                         in_data[792],
                         in_data[384],
                         in_data[591]
                    }),
            .out_data(lut_63_out)
        );

reg   lut_63_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_63_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_63_ff <= lut_63_out;
    end
end

assign out_data[63] = lut_63_ff;




// LUT : 64

wire lut_64_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110011111111111111111110111100011111111111110101111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_64
        (
            .in_data({
                         in_data[904],
                         in_data[448],
                         in_data[457],
                         in_data[989],
                         in_data[619],
                         in_data[985]
                    }),
            .out_data(lut_64_out)
        );

reg   lut_64_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_64_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_64_ff <= lut_64_out;
    end
end

assign out_data[64] = lut_64_ff;




// LUT : 65

wire lut_65_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000000000000000000000000000000100010000010100010101000000010),
            .DEVICE(DEVICE)
        )
    i_lut_65
        (
            .in_data({
                         in_data[185],
                         in_data[200],
                         in_data[21],
                         in_data[499],
                         in_data[162],
                         in_data[249]
                    }),
            .out_data(lut_65_out)
        );

reg   lut_65_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_65_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_65_ff <= lut_65_out;
    end
end

assign out_data[65] = lut_65_ff;




// LUT : 66

wire lut_66_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000001110001000100000000010001101000000001010101000000000),
            .DEVICE(DEVICE)
        )
    i_lut_66
        (
            .in_data({
                         in_data[13],
                         in_data[573],
                         in_data[921],
                         in_data[122],
                         in_data[568],
                         in_data[765]
                    }),
            .out_data(lut_66_out)
        );

reg   lut_66_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_66_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_66_ff <= lut_66_out;
    end
end

assign out_data[66] = lut_66_ff;




// LUT : 67

wire lut_67_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111100010011101111110001111101011111000110111101111100011011),
            .DEVICE(DEVICE)
        )
    i_lut_67
        (
            .in_data({
                         in_data[891],
                         in_data[391],
                         in_data[410],
                         in_data[28],
                         in_data[897],
                         in_data[695]
                    }),
            .out_data(lut_67_out)
        );

reg   lut_67_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_67_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_67_ff <= lut_67_out;
    end
end

assign out_data[67] = lut_67_ff;




// LUT : 68

wire lut_68_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000111010000000000001110010111111101000000100010010010000001),
            .DEVICE(DEVICE)
        )
    i_lut_68
        (
            .in_data({
                         in_data[903],
                         in_data[1016],
                         in_data[109],
                         in_data[516],
                         in_data[260],
                         in_data[67]
                    }),
            .out_data(lut_68_out)
        );

reg   lut_68_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_68_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_68_ff <= lut_68_out;
    end
end

assign out_data[68] = lut_68_ff;




// LUT : 69

wire lut_69_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000000000000100000000000000000000000000000000000010000000000),
            .DEVICE(DEVICE)
        )
    i_lut_69
        (
            .in_data({
                         in_data[911],
                         in_data[709],
                         in_data[441],
                         in_data[309],
                         in_data[284],
                         in_data[206]
                    }),
            .out_data(lut_69_out)
        );

reg   lut_69_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_69_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_69_ff <= lut_69_out;
    end
end

assign out_data[69] = lut_69_ff;




// LUT : 70

wire lut_70_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000010000000100000000000000001000000010001001101010001010000),
            .DEVICE(DEVICE)
        )
    i_lut_70
        (
            .in_data({
                         in_data[658],
                         in_data[582],
                         in_data[581],
                         in_data[327],
                         in_data[439],
                         in_data[280]
                    }),
            .out_data(lut_70_out)
        );

reg   lut_70_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_70_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_70_ff <= lut_70_out;
    end
end

assign out_data[70] = lut_70_ff;




// LUT : 71

wire lut_71_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001101110011000100110111011101110101011101110110011101110111),
            .DEVICE(DEVICE)
        )
    i_lut_71
        (
            .in_data({
                         in_data[623],
                         in_data[988],
                         in_data[530],
                         in_data[764],
                         in_data[732],
                         in_data[758]
                    }),
            .out_data(lut_71_out)
        );

reg   lut_71_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_71_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_71_ff <= lut_71_out;
    end
end

assign out_data[71] = lut_71_ff;




// LUT : 72

wire lut_72_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101011111111001100000111010000010000111111001111000011110100),
            .DEVICE(DEVICE)
        )
    i_lut_72
        (
            .in_data({
                         in_data[536],
                         in_data[975],
                         in_data[507],
                         in_data[324],
                         in_data[484],
                         in_data[86]
                    }),
            .out_data(lut_72_out)
        );

reg   lut_72_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_72_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_72_ff <= lut_72_out;
    end
end

assign out_data[72] = lut_72_ff;




// LUT : 73

wire lut_73_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101011111001101000101111010110101010010101001110111101011101),
            .DEVICE(DEVICE)
        )
    i_lut_73
        (
            .in_data({
                         in_data[82],
                         in_data[868],
                         in_data[234],
                         in_data[105],
                         in_data[246],
                         in_data[776]
                    }),
            .out_data(lut_73_out)
        );

reg   lut_73_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_73_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_73_ff <= lut_73_out;
    end
end

assign out_data[73] = lut_73_ff;




// LUT : 74

wire lut_74_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110011101110111011001100110000001100110010000000010001001100),
            .DEVICE(DEVICE)
        )
    i_lut_74
        (
            .in_data({
                         in_data[583],
                         in_data[254],
                         in_data[335],
                         in_data[317],
                         in_data[1008],
                         in_data[702]
                    }),
            .out_data(lut_74_out)
        );

reg   lut_74_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_74_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_74_ff <= lut_74_out;
    end
end

assign out_data[74] = lut_74_ff;




// LUT : 75

wire lut_75_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111111100110101001110001011111101111111010101111011101110111),
            .DEVICE(DEVICE)
        )
    i_lut_75
        (
            .in_data({
                         in_data[854],
                         in_data[440],
                         in_data[256],
                         in_data[775],
                         in_data[59],
                         in_data[0]
                    }),
            .out_data(lut_75_out)
        );

reg   lut_75_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_75_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_75_ff <= lut_75_out;
    end
end

assign out_data[75] = lut_75_ff;




// LUT : 76

wire lut_76_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001011110101001100111111000100110010111111000010000011001101),
            .DEVICE(DEVICE)
        )
    i_lut_76
        (
            .in_data({
                         in_data[610],
                         in_data[401],
                         in_data[69],
                         in_data[358],
                         in_data[639],
                         in_data[406]
                    }),
            .out_data(lut_76_out)
        );

reg   lut_76_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_76_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_76_ff <= lut_76_out;
    end
end

assign out_data[76] = lut_76_ff;




// LUT : 77

wire lut_77_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100010011101110000000000110101010101000101010100000000010101010),
            .DEVICE(DEVICE)
        )
    i_lut_77
        (
            .in_data({
                         in_data[196],
                         in_data[281],
                         in_data[62],
                         in_data[673],
                         in_data[325],
                         in_data[739]
                    }),
            .out_data(lut_77_out)
        );

reg   lut_77_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_77_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_77_ff <= lut_77_out;
    end
end

assign out_data[77] = lut_77_ff;




// LUT : 78

wire lut_78_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111101111111000001110000000110000111010001010110000101000101),
            .DEVICE(DEVICE)
        )
    i_lut_78
        (
            .in_data({
                         in_data[823],
                         in_data[918],
                         in_data[579],
                         in_data[369],
                         in_data[405],
                         in_data[794]
                    }),
            .out_data(lut_78_out)
        );

reg   lut_78_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_78_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_78_ff <= lut_78_out;
    end
end

assign out_data[78] = lut_78_ff;




// LUT : 79

wire lut_79_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001000000011100000101000011110000011100001111000001010000),
            .DEVICE(DEVICE)
        )
    i_lut_79
        (
            .in_data({
                         in_data[212],
                         in_data[593],
                         in_data[492],
                         in_data[865],
                         in_data[720],
                         in_data[180]
                    }),
            .out_data(lut_79_out)
        );

reg   lut_79_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_79_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_79_ff <= lut_79_out;
    end
end

assign out_data[79] = lut_79_ff;




// LUT : 80

wire lut_80_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001100000001110000111000001100110000100000011000000010000000),
            .DEVICE(DEVICE)
        )
    i_lut_80
        (
            .in_data({
                         in_data[520],
                         in_data[941],
                         in_data[670],
                         in_data[381],
                         in_data[773],
                         in_data[387]
                    }),
            .out_data(lut_80_out)
        );

reg   lut_80_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_80_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_80_ff <= lut_80_out;
    end
end

assign out_data[80] = lut_80_ff;




// LUT : 81

wire lut_81_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110011011101111101101101010111001000010110011101110001010001),
            .DEVICE(DEVICE)
        )
    i_lut_81
        (
            .in_data({
                         in_data[183],
                         in_data[710],
                         in_data[49],
                         in_data[390],
                         in_data[108],
                         in_data[584]
                    }),
            .out_data(lut_81_out)
        );

reg   lut_81_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_81_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_81_ff <= lut_81_out;
    end
end

assign out_data[81] = lut_81_ff;




// LUT : 82

wire lut_82_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011110011111111110111101100110000100000001100110001000000110001),
            .DEVICE(DEVICE)
        )
    i_lut_82
        (
            .in_data({
                         in_data[962],
                         in_data[514],
                         in_data[11],
                         in_data[453],
                         in_data[693],
                         in_data[864]
                    }),
            .out_data(lut_82_out)
        );

reg   lut_82_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_82_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_82_ff <= lut_82_out;
    end
end

assign out_data[82] = lut_82_ff;




// LUT : 83

wire lut_83_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101000011101001000001100101100010100000000000001100001010100),
            .DEVICE(DEVICE)
        )
    i_lut_83
        (
            .in_data({
                         in_data[647],
                         in_data[733],
                         in_data[178],
                         in_data[1007],
                         in_data[293],
                         in_data[714]
                    }),
            .out_data(lut_83_out)
        );

reg   lut_83_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_83_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_83_ff <= lut_83_out;
    end
end

assign out_data[83] = lut_83_ff;




// LUT : 84

wire lut_84_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010011000000100000011110000110000101010000010001100110010001100),
            .DEVICE(DEVICE)
        )
    i_lut_84
        (
            .in_data({
                         in_data[721],
                         in_data[592],
                         in_data[311],
                         in_data[442],
                         in_data[93],
                         in_data[518]
                    }),
            .out_data(lut_84_out)
        );

reg   lut_84_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_84_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_84_ff <= lut_84_out;
    end
end

assign out_data[84] = lut_84_ff;




// LUT : 85

wire lut_85_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111111111111011111101011111011111111111),
            .DEVICE(DEVICE)
        )
    i_lut_85
        (
            .in_data({
                         in_data[4],
                         in_data[386],
                         in_data[181],
                         in_data[523],
                         in_data[900],
                         in_data[270]
                    }),
            .out_data(lut_85_out)
        );

reg   lut_85_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_85_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_85_ff <= lut_85_out;
    end
end

assign out_data[85] = lut_85_ff;




// LUT : 86

wire lut_86_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111101010100111111110111111111111111000000001111111111110101),
            .DEVICE(DEVICE)
        )
    i_lut_86
        (
            .in_data({
                         in_data[398],
                         in_data[272],
                         in_data[977],
                         in_data[535],
                         in_data[68],
                         in_data[351]
                    }),
            .out_data(lut_86_out)
        );

reg   lut_86_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_86_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_86_ff <= lut_86_out;
    end
end

assign out_data[86] = lut_86_ff;




// LUT : 87

wire lut_87_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011100111111011101110001111111111111001111111111111101111111),
            .DEVICE(DEVICE)
        )
    i_lut_87
        (
            .in_data({
                         in_data[713],
                         in_data[392],
                         in_data[859],
                         in_data[819],
                         in_data[371],
                         in_data[37]
                    }),
            .out_data(lut_87_out)
        );

reg   lut_87_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_87_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_87_ff <= lut_87_out;
    end
end

assign out_data[87] = lut_87_ff;




// LUT : 88

wire lut_88_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001111100111100000010000000111000000111101011101010111110001),
            .DEVICE(DEVICE)
        )
    i_lut_88
        (
            .in_data({
                         in_data[841],
                         in_data[984],
                         in_data[607],
                         in_data[910],
                         in_data[754],
                         in_data[283]
                    }),
            .out_data(lut_88_out)
        );

reg   lut_88_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_88_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_88_ff <= lut_88_out;
    end
end

assign out_data[88] = lut_88_ff;




// LUT : 89

wire lut_89_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000100000001100100011001110111111001100100011001100110011101100),
            .DEVICE(DEVICE)
        )
    i_lut_89
        (
            .in_data({
                         in_data[1005],
                         in_data[969],
                         in_data[837],
                         in_data[945],
                         in_data[1002],
                         in_data[624]
                    }),
            .out_data(lut_89_out)
        );

reg   lut_89_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_89_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_89_ff <= lut_89_out;
    end
end

assign out_data[89] = lut_89_ff;




// LUT : 90

wire lut_90_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100011011111111101010111000110111101111111111011001111111111100),
            .DEVICE(DEVICE)
        )
    i_lut_90
        (
            .in_data({
                         in_data[266],
                         in_data[839],
                         in_data[239],
                         in_data[295],
                         in_data[377],
                         in_data[981]
                    }),
            .out_data(lut_90_out)
        );

reg   lut_90_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_90_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_90_ff <= lut_90_out;
    end
end

assign out_data[90] = lut_90_ff;




// LUT : 91

wire lut_91_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111110001001100110011111111111111111101010111111101),
            .DEVICE(DEVICE)
        )
    i_lut_91
        (
            .in_data({
                         in_data[802],
                         in_data[231],
                         in_data[980],
                         in_data[596],
                         in_data[942],
                         in_data[417]
                    }),
            .out_data(lut_91_out)
        );

reg   lut_91_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_91_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_91_ff <= lut_91_out;
    end
end

assign out_data[91] = lut_91_ff;




// LUT : 92

wire lut_92_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110001111110110110000011011111010010111010101111100000000),
            .DEVICE(DEVICE)
        )
    i_lut_92
        (
            .in_data({
                         in_data[1],
                         in_data[61],
                         in_data[952],
                         in_data[508],
                         in_data[808],
                         in_data[810]
                    }),
            .out_data(lut_92_out)
        );

reg   lut_92_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_92_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_92_ff <= lut_92_out;
    end
end

assign out_data[92] = lut_92_ff;




// LUT : 93

wire lut_93_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001000100011000001110000001100000011111110100000000000000010),
            .DEVICE(DEVICE)
        )
    i_lut_93
        (
            .in_data({
                         in_data[795],
                         in_data[960],
                         in_data[876],
                         in_data[471],
                         in_data[226],
                         in_data[110]
                    }),
            .out_data(lut_93_out)
        );

reg   lut_93_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_93_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_93_ff <= lut_93_out;
    end
end

assign out_data[93] = lut_93_ff;




// LUT : 94

wire lut_94_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100010001101000010100001011000001111100110110011101100011000),
            .DEVICE(DEVICE)
        )
    i_lut_94
        (
            .in_data({
                         in_data[889],
                         in_data[341],
                         in_data[781],
                         in_data[143],
                         in_data[616],
                         in_data[554]
                    }),
            .out_data(lut_94_out)
        );

reg   lut_94_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_94_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_94_ff <= lut_94_out;
    end
end

assign out_data[94] = lut_94_ff;




// LUT : 95

wire lut_95_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010011110011110010011101111101111101100001010101011001011010),
            .DEVICE(DEVICE)
        )
    i_lut_95
        (
            .in_data({
                         in_data[679],
                         in_data[731],
                         in_data[986],
                         in_data[997],
                         in_data[449],
                         in_data[456]
                    }),
            .out_data(lut_95_out)
        );

reg   lut_95_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_95_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_95_ff <= lut_95_out;
    end
end

assign out_data[95] = lut_95_ff;




// LUT : 96

wire lut_96_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001000000000100011111000100000000000000000000000110000000000),
            .DEVICE(DEVICE)
        )
    i_lut_96
        (
            .in_data({
                         in_data[552],
                         in_data[347],
                         in_data[32],
                         in_data[150],
                         in_data[632],
                         in_data[321]
                    }),
            .out_data(lut_96_out)
        );

reg   lut_96_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_96_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_96_ff <= lut_96_out;
    end
end

assign out_data[96] = lut_96_ff;




// LUT : 97

wire lut_97_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101011000100111111101111111111111110110111011111110111111111),
            .DEVICE(DEVICE)
        )
    i_lut_97
        (
            .in_data({
                         in_data[416],
                         in_data[279],
                         in_data[378],
                         in_data[495],
                         in_data[762],
                         in_data[828]
                    }),
            .out_data(lut_97_out)
        );

reg   lut_97_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_97_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_97_ff <= lut_97_out;
    end
end

assign out_data[97] = lut_97_ff;




// LUT : 98

wire lut_98_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000011011000010111011101110101010000010101010001010100010101),
            .DEVICE(DEVICE)
        )
    i_lut_98
        (
            .in_data({
                         in_data[362],
                         in_data[614],
                         in_data[524],
                         in_data[314],
                         in_data[219],
                         in_data[71]
                    }),
            .out_data(lut_98_out)
        );

reg   lut_98_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_98_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_98_ff <= lut_98_out;
    end
end

assign out_data[98] = lut_98_ff;




// LUT : 99

wire lut_99_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101010101010000010000010111101000000000010100000000000001111),
            .DEVICE(DEVICE)
        )
    i_lut_99
        (
            .in_data({
                         in_data[948],
                         in_data[763],
                         in_data[51],
                         in_data[838],
                         in_data[156],
                         in_data[75]
                    }),
            .out_data(lut_99_out)
        );

reg   lut_99_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_99_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_99_ff <= lut_99_out;
    end
end

assign out_data[99] = lut_99_ff;




// LUT : 100

wire lut_100_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110011001100100101110110110111000000110000001010000101111100),
            .DEVICE(DEVICE)
        )
    i_lut_100
        (
            .in_data({
                         in_data[74],
                         in_data[385],
                         in_data[821],
                         in_data[697],
                         in_data[906],
                         in_data[567]
                    }),
            .out_data(lut_100_out)
        );

reg   lut_100_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_100_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_100_ff <= lut_100_out;
    end
end

assign out_data[100] = lut_100_ff;




// LUT : 101

wire lut_101_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001011111111001100111111111110111011111111110010001010101011),
            .DEVICE(DEVICE)
        )
    i_lut_101
        (
            .in_data({
                         in_data[46],
                         in_data[103],
                         in_data[698],
                         in_data[135],
                         in_data[8],
                         in_data[621]
                    }),
            .out_data(lut_101_out)
        );

reg   lut_101_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_101_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_101_ff <= lut_101_out;
    end
end

assign out_data[101] = lut_101_ff;




// LUT : 102

wire lut_102_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001001100011011000101110001111100000011000000110000000100000000),
            .DEVICE(DEVICE)
        )
    i_lut_102
        (
            .in_data({
                         in_data[824],
                         in_data[668],
                         in_data[641],
                         in_data[479],
                         in_data[769],
                         in_data[835]
                    }),
            .out_data(lut_102_out)
        );

reg   lut_102_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_102_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_102_ff <= lut_102_out;
    end
end

assign out_data[102] = lut_102_ff;




// LUT : 103

wire lut_103_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001011101011111011111100111111111000110110101101111011111110),
            .DEVICE(DEVICE)
        )
    i_lut_103
        (
            .in_data({
                         in_data[675],
                         in_data[618],
                         in_data[120],
                         in_data[588],
                         in_data[800],
                         in_data[885]
                    }),
            .out_data(lut_103_out)
        );

reg   lut_103_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_103_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_103_ff <= lut_103_out;
    end
end

assign out_data[103] = lut_103_ff;




// LUT : 104

wire lut_104_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011111111111111111111111111111110101111101011111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_104
        (
            .in_data({
                         in_data[235],
                         in_data[52],
                         in_data[411],
                         in_data[558],
                         in_data[287],
                         in_data[140]
                    }),
            .out_data(lut_104_out)
        );

reg   lut_104_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_104_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_104_ff <= lut_104_out;
    end
end

assign out_data[104] = lut_104_ff;




// LUT : 105

wire lut_105_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111010111011011111111111101011111110111),
            .DEVICE(DEVICE)
        )
    i_lut_105
        (
            .in_data({
                         in_data[496],
                         in_data[244],
                         in_data[715],
                         in_data[553],
                         in_data[127],
                         in_data[194]
                    }),
            .out_data(lut_105_out)
        );

reg   lut_105_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_105_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_105_ff <= lut_105_out;
    end
end

assign out_data[105] = lut_105_ff;




// LUT : 106

wire lut_106_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100010000000100000001100000000000000101000101010100011010000),
            .DEVICE(DEVICE)
        )
    i_lut_106
        (
            .in_data({
                         in_data[515],
                         in_data[737],
                         in_data[915],
                         in_data[87],
                         in_data[929],
                         in_data[893]
                    }),
            .out_data(lut_106_out)
        );

reg   lut_106_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_106_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_106_ff <= lut_106_out;
    end
end

assign out_data[106] = lut_106_ff;




// LUT : 107

wire lut_107_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000100010000100000000001001000000111001010001100110000000000),
            .DEVICE(DEVICE)
        )
    i_lut_107
        (
            .in_data({
                         in_data[853],
                         in_data[768],
                         in_data[188],
                         in_data[498],
                         in_data[772],
                         in_data[240]
                    }),
            .out_data(lut_107_out)
        );

reg   lut_107_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_107_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_107_ff <= lut_107_out;
    end
end

assign out_data[107] = lut_107_ff;




// LUT : 108

wire lut_108_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010100010001000100000000000001110101011101110111010100110001),
            .DEVICE(DEVICE)
        )
    i_lut_108
        (
            .in_data({
                         in_data[569],
                         in_data[716],
                         in_data[944],
                         in_data[476],
                         in_data[1003],
                         in_data[202]
                    }),
            .out_data(lut_108_out)
        );

reg   lut_108_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_108_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_108_ff <= lut_108_out;
    end
end

assign out_data[108] = lut_108_ff;




// LUT : 109

wire lut_109_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110101010101110111111101111101000100010001001101111011111110),
            .DEVICE(DEVICE)
        )
    i_lut_109
        (
            .in_data({
                         in_data[722],
                         in_data[917],
                         in_data[556],
                         in_data[36],
                         in_data[72],
                         in_data[115]
                    }),
            .out_data(lut_109_out)
        );

reg   lut_109_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_109_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_109_ff <= lut_109_out;
    end
end

assign out_data[109] = lut_109_ff;




// LUT : 110

wire lut_110_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010101000000010000000100000001000101000000001100000001100000),
            .DEVICE(DEVICE)
        )
    i_lut_110
        (
            .in_data({
                         in_data[469],
                         in_data[734],
                         in_data[884],
                         in_data[955],
                         in_data[438],
                         in_data[273]
                    }),
            .out_data(lut_110_out)
        );

reg   lut_110_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_110_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_110_ff <= lut_110_out;
    end
end

assign out_data[110] = lut_110_ff;




// LUT : 111

wire lut_111_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111101010111010111000101000001110111000000101111100100101000),
            .DEVICE(DEVICE)
        )
    i_lut_111
        (
            .in_data({
                         in_data[308],
                         in_data[124],
                         in_data[259],
                         in_data[315],
                         in_data[430],
                         in_data[253]
                    }),
            .out_data(lut_111_out)
        );

reg   lut_111_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_111_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_111_ff <= lut_111_out;
    end
end

assign out_data[111] = lut_111_ff;




// LUT : 112

wire lut_112_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000000100000011100111111001101000100111101000111000011110000),
            .DEVICE(DEVICE)
        )
    i_lut_112
        (
            .in_data({
                         in_data[278],
                         in_data[660],
                         in_data[798],
                         in_data[121],
                         in_data[615],
                         in_data[831]
                    }),
            .out_data(lut_112_out)
        );

reg   lut_112_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_112_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_112_ff <= lut_112_out;
    end
end

assign out_data[112] = lut_112_ff;




// LUT : 113

wire lut_113_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110011111111010101000101010011111000000110000001000100010001),
            .DEVICE(DEVICE)
        )
    i_lut_113
        (
            .in_data({
                         in_data[493],
                         in_data[881],
                         in_data[81],
                         in_data[1000],
                         in_data[157],
                         in_data[80]
                    }),
            .out_data(lut_113_out)
        );

reg   lut_113_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_113_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_113_ff <= lut_113_out;
    end
end

assign out_data[113] = lut_113_ff;




// LUT : 114

wire lut_114_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101111101110111111111111111100000000110111001010111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_114
        (
            .in_data({
                         in_data[224],
                         in_data[78],
                         in_data[248],
                         in_data[230],
                         in_data[968],
                         in_data[153]
                    }),
            .out_data(lut_114_out)
        );

reg   lut_114_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_114_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_114_ff <= lut_114_out;
    end
end

assign out_data[114] = lut_114_ff;




// LUT : 115

wire lut_115_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000011000100110101001101010000000000000000000100000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_115
        (
            .in_data({
                         in_data[198],
                         in_data[752],
                         in_data[258],
                         in_data[10],
                         in_data[1014],
                         in_data[376]
                    }),
            .out_data(lut_115_out)
        );

reg   lut_115_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_115_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_115_ff <= lut_115_out;
    end
end

assign out_data[115] = lut_115_ff;




// LUT : 116

wire lut_116_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101100101001101010110010110010101010000010100000000000000011),
            .DEVICE(DEVICE)
        )
    i_lut_116
        (
            .in_data({
                         in_data[112],
                         in_data[27],
                         in_data[30],
                         in_data[559],
                         in_data[685],
                         in_data[275]
                    }),
            .out_data(lut_116_out)
        );

reg   lut_116_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_116_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_116_ff <= lut_116_out;
    end
end

assign out_data[116] = lut_116_ff;




// LUT : 117

wire lut_117_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000110010000100100010101000000000000000000001010100001011),
            .DEVICE(DEVICE)
        )
    i_lut_117
        (
            .in_data({
                         in_data[546],
                         in_data[760],
                         in_data[847],
                         in_data[799],
                         in_data[594],
                         in_data[1017]
                    }),
            .out_data(lut_117_out)
        );

reg   lut_117_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_117_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_117_ff <= lut_117_out;
    end
end

assign out_data[117] = lut_117_ff;




// LUT : 118

wire lut_118_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000010001010000010101001000010001001100110101000101),
            .DEVICE(DEVICE)
        )
    i_lut_118
        (
            .in_data({
                         in_data[612],
                         in_data[790],
                         in_data[780],
                         in_data[274],
                         in_data[177],
                         in_data[182]
                    }),
            .out_data(lut_118_out)
        );

reg   lut_118_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_118_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_118_ff <= lut_118_out;
    end
end

assign out_data[118] = lut_118_ff;




// LUT : 119

wire lut_119_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111101000111111110011010001001111111101000100110100111000),
            .DEVICE(DEVICE)
        )
    i_lut_119
        (
            .in_data({
                         in_data[645],
                         in_data[974],
                         in_data[412],
                         in_data[700],
                         in_data[285],
                         in_data[861]
                    }),
            .out_data(lut_119_out)
        );

reg   lut_119_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_119_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_119_ff <= lut_119_out;
    end
end

assign out_data[119] = lut_119_ff;




// LUT : 120

wire lut_120_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000111111100111111111111111100000000110011100000000111001111),
            .DEVICE(DEVICE)
        )
    i_lut_120
        (
            .in_data({
                         in_data[425],
                         in_data[241],
                         in_data[743],
                         in_data[205],
                         in_data[383],
                         in_data[9]
                    }),
            .out_data(lut_120_out)
        );

reg   lut_120_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_120_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_120_ff <= lut_120_out;
    end
end

assign out_data[120] = lut_120_ff;




// LUT : 121

wire lut_121_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111111111111100111011101111110011101110),
            .DEVICE(DEVICE)
        )
    i_lut_121
        (
            .in_data({
                         in_data[644],
                         in_data[866],
                         in_data[38],
                         in_data[843],
                         in_data[676],
                         in_data[862]
                    }),
            .out_data(lut_121_out)
        );

reg   lut_121_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_121_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_121_ff <= lut_121_out;
    end
end

assign out_data[121] = lut_121_ff;




// LUT : 122

wire lut_122_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111100010001000010110001000100000001000100010000000100010001),
            .DEVICE(DEVICE)
        )
    i_lut_122
        (
            .in_data({
                         in_data[1012],
                         in_data[643],
                         in_data[264],
                         in_data[503],
                         in_data[807],
                         in_data[872]
                    }),
            .out_data(lut_122_out)
        );

reg   lut_122_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_122_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_122_ff <= lut_122_out;
    end
end

assign out_data[122] = lut_122_ff;




// LUT : 123

wire lut_123_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111011111111000010100100111000000000000000000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_123
        (
            .in_data({
                         in_data[712],
                         in_data[669],
                         in_data[329],
                         in_data[199],
                         in_data[468],
                         in_data[708]
                    }),
            .out_data(lut_123_out)
        );

reg   lut_123_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_123_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_123_ff <= lut_123_out;
    end
end

assign out_data[123] = lut_123_ff;




// LUT : 124

wire lut_124_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001011111101111111111111110100111011001111111000111011111000),
            .DEVICE(DEVICE)
        )
    i_lut_124
        (
            .in_data({
                         in_data[319],
                         in_data[312],
                         in_data[145],
                         in_data[683],
                         in_data[477],
                         in_data[354]
                    }),
            .out_data(lut_124_out)
        );

reg   lut_124_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_124_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_124_ff <= lut_124_out;
    end
end

assign out_data[124] = lut_124_ff;




// LUT : 125

wire lut_125_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000101101000000001100111100100011001100110000000100010001),
            .DEVICE(DEVICE)
        )
    i_lut_125
        (
            .in_data({
                         in_data[555],
                         in_data[344],
                         in_data[656],
                         in_data[998],
                         in_data[1004],
                         in_data[250]
                    }),
            .out_data(lut_125_out)
        );

reg   lut_125_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_125_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_125_ff <= lut_125_out;
    end
end

assign out_data[125] = lut_125_ff;




// LUT : 126

wire lut_126_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110011100010000100001010001100010000000111010101000010001100),
            .DEVICE(DEVICE)
        )
    i_lut_126
        (
            .in_data({
                         in_data[47],
                         in_data[735],
                         in_data[661],
                         in_data[711],
                         in_data[24],
                         in_data[197]
                    }),
            .out_data(lut_126_out)
        );

reg   lut_126_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_126_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_126_ff <= lut_126_out;
    end
end

assign out_data[126] = lut_126_ff;




// LUT : 127

wire lut_127_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001011101110111001100110000101100001010001010110000001000101011),
            .DEVICE(DEVICE)
        )
    i_lut_127
        (
            .in_data({
                         in_data[263],
                         in_data[159],
                         in_data[613],
                         in_data[901],
                         in_data[855],
                         in_data[625]
                    }),
            .out_data(lut_127_out)
        );

reg   lut_127_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_127_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_127_ff <= lut_127_out;
    end
end

assign out_data[127] = lut_127_ff;




// LUT : 128

wire lut_128_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000011000000110001000000000001000100010000000100010111100101111),
            .DEVICE(DEVICE)
        )
    i_lut_128
        (
            .in_data({
                         in_data[34],
                         in_data[443],
                         in_data[525],
                         in_data[631],
                         in_data[407],
                         in_data[356]
                    }),
            .out_data(lut_128_out)
        );

reg   lut_128_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_128_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_128_ff <= lut_128_out;
    end
end

assign out_data[128] = lut_128_ff;




// LUT : 129

wire lut_129_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111010010100101111100001011101111110000000000111011),
            .DEVICE(DEVICE)
        )
    i_lut_129
        (
            .in_data({
                         in_data[189],
                         in_data[88],
                         in_data[348],
                         in_data[730],
                         in_data[517],
                         in_data[346]
                    }),
            .out_data(lut_129_out)
        );

reg   lut_129_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_129_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_129_ff <= lut_129_out;
    end
end

assign out_data[129] = lut_129_ff;




// LUT : 130

wire lut_130_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011111110111111100011111011101110011111101110111000001110011),
            .DEVICE(DEVICE)
        )
    i_lut_130
        (
            .in_data({
                         in_data[220],
                         in_data[748],
                         in_data[659],
                         in_data[16],
                         in_data[144],
                         in_data[766]
                    }),
            .out_data(lut_130_out)
        );

reg   lut_130_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_130_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_130_ff <= lut_130_out;
    end
end

assign out_data[130] = lut_130_ff;




// LUT : 131

wire lut_131_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111100000000111111111010111111001110111111001001101011101010),
            .DEVICE(DEVICE)
        )
    i_lut_131
        (
            .in_data({
                         in_data[292],
                         in_data[877],
                         in_data[470],
                         in_data[931],
                         in_data[396],
                         in_data[42]
                    }),
            .out_data(lut_131_out)
        );

reg   lut_131_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_131_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_131_ff <= lut_131_out;
    end
end

assign out_data[131] = lut_131_ff;




// LUT : 132

wire lut_132_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110011000100000101001110110100110000010011100011001000110111),
            .DEVICE(DEVICE)
        )
    i_lut_132
        (
            .in_data({
                         in_data[992],
                         in_data[727],
                         in_data[55],
                         in_data[12],
                         in_data[164],
                         in_data[175]
                    }),
            .out_data(lut_132_out)
        );

reg   lut_132_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_132_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_132_ff <= lut_132_out;
    end
end

assign out_data[132] = lut_132_ff;




// LUT : 133

wire lut_133_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000011101000111010001110111111111000111011101110100011001010),
            .DEVICE(DEVICE)
        )
    i_lut_133
        (
            .in_data({
                         in_data[316],
                         in_data[301],
                         in_data[538],
                         in_data[363],
                         in_data[723],
                         in_data[118]
                    }),
            .out_data(lut_133_out)
        );

reg   lut_133_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_133_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_133_ff <= lut_133_out;
    end
end

assign out_data[133] = lut_133_ff;




// LUT : 134

wire lut_134_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110001111110111000001100011111101110011111101110011011000),
            .DEVICE(DEVICE)
        )
    i_lut_134
        (
            .in_data({
                         in_data[413],
                         in_data[41],
                         in_data[813],
                         in_data[869],
                         in_data[216],
                         in_data[875]
                    }),
            .out_data(lut_134_out)
        );

reg   lut_134_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_134_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_134_ff <= lut_134_out;
    end
end

assign out_data[134] = lut_134_ff;




// LUT : 135

wire lut_135_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000010011000100111000011111001000000100000000000000001110000),
            .DEVICE(DEVICE)
        )
    i_lut_135
        (
            .in_data({
                         in_data[626],
                         in_data[215],
                         in_data[599],
                         in_data[73],
                         in_data[500],
                         in_data[342]
                    }),
            .out_data(lut_135_out)
        );

reg   lut_135_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_135_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_135_ff <= lut_135_out;
    end
end

assign out_data[135] = lut_135_ff;




// LUT : 136

wire lut_136_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100000000100101011111011111111111110111111111111111111101111),
            .DEVICE(DEVICE)
        )
    i_lut_136
        (
            .in_data({
                         in_data[562],
                         in_data[825],
                         in_data[575],
                         in_data[119],
                         in_data[718],
                         in_data[445]
                    }),
            .out_data(lut_136_out)
        );

reg   lut_136_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_136_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_136_ff <= lut_136_out;
    end
end

assign out_data[136] = lut_136_ff;




// LUT : 137

wire lut_137_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111101001101100010111011010100110111111011110001100100111011),
            .DEVICE(DEVICE)
        )
    i_lut_137
        (
            .in_data({
                         in_data[245],
                         in_data[426],
                         in_data[826],
                         in_data[845],
                         in_data[225],
                         in_data[534]
                    }),
            .out_data(lut_137_out)
        );

reg   lut_137_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_137_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_137_ff <= lut_137_out;
    end
end

assign out_data[137] = lut_137_ff;




// LUT : 138

wire lut_138_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000011001100110011001110100101000000110011111100100111010101),
            .DEVICE(DEVICE)
        )
    i_lut_138
        (
            .in_data({
                         in_data[5],
                         in_data[191],
                         in_data[90],
                         in_data[848],
                         in_data[265],
                         in_data[657]
                    }),
            .out_data(lut_138_out)
        );

reg   lut_138_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_138_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_138_ff <= lut_138_out;
    end
end

assign out_data[138] = lut_138_ff;




// LUT : 139

wire lut_139_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101101111111110000110111111111100011000011110101010111100111111),
            .DEVICE(DEVICE)
        )
    i_lut_139
        (
            .in_data({
                         in_data[1019],
                         in_data[755],
                         in_data[815],
                         in_data[630],
                         in_data[682],
                         in_data[842]
                    }),
            .out_data(lut_139_out)
        );

reg   lut_139_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_139_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_139_ff <= lut_139_out;
    end
end

assign out_data[139] = lut_139_ff;




// LUT : 140

wire lut_140_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111110111101101111111001110111111101111111011011100111011101),
            .DEVICE(DEVICE)
        )
    i_lut_140
        (
            .in_data({
                         in_data[979],
                         in_data[104],
                         in_data[464],
                         in_data[91],
                         in_data[343],
                         in_data[767]
                    }),
            .out_data(lut_140_out)
        );

reg   lut_140_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_140_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_140_ff <= lut_140_out;
    end
end

assign out_data[140] = lut_140_ff;




// LUT : 141

wire lut_141_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111000000000111011101000011011000100000000000110001000000000),
            .DEVICE(DEVICE)
        )
    i_lut_141
        (
            .in_data({
                         in_data[429],
                         in_data[483],
                         in_data[474],
                         in_data[597],
                         in_data[550],
                         in_data[305]
                    }),
            .out_data(lut_141_out)
        );

reg   lut_141_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_141_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_141_ff <= lut_141_out;
    end
end

assign out_data[141] = lut_141_ff;




// LUT : 142

wire lut_142_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111011111110011111001111111111110111111101011111100111111101),
            .DEVICE(DEVICE)
        )
    i_lut_142
        (
            .in_data({
                         in_data[40],
                         in_data[664],
                         in_data[505],
                         in_data[201],
                         in_data[50],
                         in_data[545]
                    }),
            .out_data(lut_142_out)
        );

reg   lut_142_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_142_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_142_ff <= lut_142_out;
    end
end

assign out_data[142] = lut_142_ff;




// LUT : 143

wire lut_143_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000011010000110000100000101111111110110110101100111111111010),
            .DEVICE(DEVICE)
        )
    i_lut_143
        (
            .in_data({
                         in_data[681],
                         in_data[880],
                         in_data[450],
                         in_data[310],
                         in_data[577],
                         in_data[380]
                    }),
            .out_data(lut_143_out)
        );

reg   lut_143_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_143_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_143_ff <= lut_143_out;
    end
end

assign out_data[143] = lut_143_ff;




// LUT : 144

wire lut_144_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110111111010111110100111111111011111100111111110100000001),
            .DEVICE(DEVICE)
        )
    i_lut_144
        (
            .in_data({
                         in_data[791],
                         in_data[991],
                         in_data[674],
                         in_data[57],
                         in_data[257],
                         in_data[829]
                    }),
            .out_data(lut_144_out)
        );

reg   lut_144_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_144_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_144_ff <= lut_144_out;
    end
end

assign out_data[144] = lut_144_ff;




// LUT : 145

wire lut_145_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111000000100010101111111111001000111010001000100010),
            .DEVICE(DEVICE)
        )
    i_lut_145
        (
            .in_data({
                         in_data[485],
                         in_data[35],
                         in_data[137],
                         in_data[784],
                         in_data[454],
                         in_data[331]
                    }),
            .out_data(lut_145_out)
        );

reg   lut_145_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_145_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_145_ff <= lut_145_out;
    end
end

assign out_data[145] = lut_145_ff;




// LUT : 146

wire lut_146_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010000010100110110110000111111010001111111111111111101111101),
            .DEVICE(DEVICE)
        )
    i_lut_146
        (
            .in_data({
                         in_data[1018],
                         in_data[366],
                         in_data[23],
                         in_data[186],
                         in_data[542],
                         in_data[218]
                    }),
            .out_data(lut_146_out)
        );

reg   lut_146_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_146_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_146_ff <= lut_146_out;
    end
end

assign out_data[146] = lut_146_ff;




// LUT : 147

wire lut_147_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111111111111111111100011111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_147
        (
            .in_data({
                         in_data[598],
                         in_data[919],
                         in_data[447],
                         in_data[133],
                         in_data[595],
                         in_data[585]
                    }),
            .out_data(lut_147_out)
        );

reg   lut_147_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_147_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_147_ff <= lut_147_out;
    end
end

assign out_data[147] = lut_147_ff;




// LUT : 148

wire lut_148_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000001001100110000001101110011000010010001001101000011000100),
            .DEVICE(DEVICE)
        )
    i_lut_148
        (
            .in_data({
                         in_data[688],
                         in_data[1015],
                         in_data[951],
                         in_data[719],
                         in_data[422],
                         in_data[261]
                    }),
            .out_data(lut_148_out)
        );

reg   lut_148_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_148_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_148_ff <= lut_148_out;
    end
end

assign out_data[148] = lut_148_ff;




// LUT : 149

wire lut_149_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111101111111011001010101010101010010010111110101000001010111),
            .DEVICE(DEVICE)
        )
    i_lut_149
        (
            .in_data({
                         in_data[409],
                         in_data[860],
                         in_data[149],
                         in_data[922],
                         in_data[940],
                         in_data[1023]
                    }),
            .out_data(lut_149_out)
        );

reg   lut_149_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_149_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_149_ff <= lut_149_out;
    end
end

assign out_data[149] = lut_149_ff;




// LUT : 150

wire lut_150_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101001101010100000010001100000001010101110100000010111111100000),
            .DEVICE(DEVICE)
        )
    i_lut_150
        (
            .in_data({
                         in_data[1001],
                         in_data[45],
                         in_data[586],
                         in_data[740],
                         in_data[927],
                         in_data[17]
                    }),
            .out_data(lut_150_out)
        );

reg   lut_150_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_150_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_150_ff <= lut_150_out;
    end
end

assign out_data[150] = lut_150_ff;




// LUT : 151

wire lut_151_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110111100101010011111100000001011011111110111111111111111011010),
            .DEVICE(DEVICE)
        )
    i_lut_151
        (
            .in_data({
                         in_data[65],
                         in_data[801],
                         in_data[187],
                         in_data[475],
                         in_data[971],
                         in_data[357]
                    }),
            .out_data(lut_151_out)
        );

reg   lut_151_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_151_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_151_ff <= lut_151_out;
    end
end

assign out_data[151] = lut_151_ff;




// LUT : 152

wire lut_152_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110011001000100000001111101000011110000000001100100000110000),
            .DEVICE(DEVICE)
        )
    i_lut_152
        (
            .in_data({
                         in_data[691],
                         in_data[814],
                         in_data[636],
                         in_data[587],
                         in_data[462],
                         in_data[204]
                    }),
            .out_data(lut_152_out)
        );

reg   lut_152_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_152_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_152_ff <= lut_152_out;
    end
end

assign out_data[152] = lut_152_ff;




// LUT : 153

wire lut_153_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111111111111101111111111111111110111111111111111010111111111),
            .DEVICE(DEVICE)
        )
    i_lut_153
        (
            .in_data({
                         in_data[176],
                         in_data[672],
                         in_data[323],
                         in_data[99],
                         in_data[816],
                         in_data[961]
                    }),
            .out_data(lut_153_out)
        );

reg   lut_153_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_153_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_153_ff <= lut_153_out;
    end
end

assign out_data[153] = lut_153_ff;




// LUT : 154

wire lut_154_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010011110110101000111010001000100011111000000100001001100000001),
            .DEVICE(DEVICE)
        )
    i_lut_154
        (
            .in_data({
                         in_data[227],
                         in_data[26],
                         in_data[48],
                         in_data[744],
                         in_data[547],
                         in_data[195]
                    }),
            .out_data(lut_154_out)
        );

reg   lut_154_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_154_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_154_ff <= lut_154_out;
    end
end

assign out_data[154] = lut_154_ff;




// LUT : 155

wire lut_155_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011101100000000000000000000000011011110111011100000000000000100),
            .DEVICE(DEVICE)
        )
    i_lut_155
        (
            .in_data({
                         in_data[446],
                         in_data[14],
                         in_data[646],
                         in_data[132],
                         in_data[489],
                         in_data[751]
                    }),
            .out_data(lut_155_out)
        );

reg   lut_155_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_155_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_155_ff <= lut_155_out;
    end
end

assign out_data[155] = lut_155_ff;




// LUT : 156

wire lut_156_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110101010101000000000000010101010101010101010000000001000101),
            .DEVICE(DEVICE)
        )
    i_lut_156
        (
            .in_data({
                         in_data[741],
                         in_data[192],
                         in_data[428],
                         in_data[15],
                         in_data[954],
                         in_data[397]
                    }),
            .out_data(lut_156_out)
        );

reg   lut_156_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_156_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_156_ff <= lut_156_out;
    end
end

assign out_data[156] = lut_156_ff;




// LUT : 157

wire lut_157_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000011001101111010111101110111001101111111111100110010010001),
            .DEVICE(DEVICE)
        )
    i_lut_157
        (
            .in_data({
                         in_data[747],
                         in_data[167],
                         in_data[3],
                         in_data[349],
                         in_data[100],
                         in_data[965]
                    }),
            .out_data(lut_157_out)
        );

reg   lut_157_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_157_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_157_ff <= lut_157_out;
    end
end

assign out_data[157] = lut_157_ff;




// LUT : 158

wire lut_158_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111111100000000101010010000101110101111),
            .DEVICE(DEVICE)
        )
    i_lut_158
        (
            .in_data({
                         in_data[909],
                         in_data[139],
                         in_data[214],
                         in_data[421],
                         in_data[705],
                         in_data[1022]
                    }),
            .out_data(lut_158_out)
        );

reg   lut_158_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_158_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_158_ff <= lut_158_out;
    end
end

assign out_data[158] = lut_158_ff;




// LUT : 159

wire lut_159_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110000100000011111111110111001011111100011100111111111111110100),
            .DEVICE(DEVICE)
        )
    i_lut_159
        (
            .in_data({
                         in_data[878],
                         in_data[207],
                         in_data[533],
                         in_data[345],
                         in_data[830],
                         in_data[551]
                    }),
            .out_data(lut_159_out)
        );

reg   lut_159_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_159_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_159_ff <= lut_159_out;
    end
end

assign out_data[159] = lut_159_ff;




// LUT : 160

wire lut_160_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000000110010000000000010000011111111001100000010001000100000),
            .DEVICE(DEVICE)
        )
    i_lut_160
        (
            .in_data({
                         in_data[908],
                         in_data[66],
                         in_data[680],
                         in_data[222],
                         in_data[653],
                         in_data[770]
                    }),
            .out_data(lut_160_out)
        );

reg   lut_160_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_160_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_160_ff <= lut_160_out;
    end
end

assign out_data[160] = lut_160_ff;




// LUT : 161

wire lut_161_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011101010101101100000011101111111111001101011011111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_161
        (
            .in_data({
                         in_data[403],
                         in_data[94],
                         in_data[251],
                         in_data[654],
                         in_data[707],
                         in_data[414]
                    }),
            .out_data(lut_161_out)
        );

reg   lut_161_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_161_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_161_ff <= lut_161_out;
    end
end

assign out_data[161] = lut_161_ff;




// LUT : 162

wire lut_162_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000010111000001100000000000000000000101110000001),
            .DEVICE(DEVICE)
        )
    i_lut_162
        (
            .in_data({
                         in_data[486],
                         in_data[994],
                         in_data[262],
                         in_data[519],
                         in_data[451],
                         in_data[355]
                    }),
            .out_data(lut_162_out)
        );

reg   lut_162_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_162_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_162_ff <= lut_162_out;
    end
end

assign out_data[162] = lut_162_ff;




// LUT : 163

wire lut_163_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011101111111010101010101010101111111011111110101110100011111),
            .DEVICE(DEVICE)
        )
    i_lut_163
        (
            .in_data({
                         in_data[753],
                         in_data[25],
                         in_data[867],
                         in_data[211],
                         in_data[541],
                         in_data[857]
                    }),
            .out_data(lut_163_out)
        );

reg   lut_163_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_163_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_163_ff <= lut_163_out;
    end
end

assign out_data[163] = lut_163_ff;




// LUT : 164

wire lut_164_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000100000000110100001100000100000001100101001111101111101111),
            .DEVICE(DEVICE)
        )
    i_lut_164
        (
            .in_data({
                         in_data[89],
                         in_data[684],
                         in_data[871],
                         in_data[289],
                         in_data[382],
                         in_data[243]
                    }),
            .out_data(lut_164_out)
        );

reg   lut_164_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_164_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_164_ff <= lut_164_out;
    end
end

assign out_data[164] = lut_164_ff;




// LUT : 165

wire lut_165_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111101111111110011010101111111111111010110101111110101011111),
            .DEVICE(DEVICE)
        )
    i_lut_165
        (
            .in_data({
                         in_data[949],
                         in_data[834],
                         in_data[19],
                         in_data[846],
                         in_data[339],
                         in_data[690]
                    }),
            .out_data(lut_165_out)
        );

reg   lut_165_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_165_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_165_ff <= lut_165_out;
    end
end

assign out_data[165] = lut_165_ff;




// LUT : 166

wire lut_166_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000100001000110110000000100010011001000110011),
            .DEVICE(DEVICE)
        )
    i_lut_166
        (
            .in_data({
                         in_data[926],
                         in_data[282],
                         in_data[978],
                         in_data[947],
                         in_data[154],
                         in_data[434]
                    }),
            .out_data(lut_166_out)
        );

reg   lut_166_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_166_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_166_ff <= lut_166_out;
    end
end

assign out_data[166] = lut_166_ff;




// LUT : 167

wire lut_167_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110111111111010011001111111100111101111111110100111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_167
        (
            .in_data({
                         in_data[379],
                         in_data[892],
                         in_data[161],
                         in_data[563],
                         in_data[532],
                         in_data[687]
                    }),
            .out_data(lut_167_out)
        );

reg   lut_167_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_167_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_167_ff <= lut_167_out;
    end
end

assign out_data[167] = lut_167_ff;




// LUT : 168

wire lut_168_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101111110011111100110111000111111111111101011111111101110001),
            .DEVICE(DEVICE)
        )
    i_lut_168
        (
            .in_data({
                         in_data[996],
                         in_data[233],
                         in_data[1011],
                         in_data[1006],
                         in_data[694],
                         in_data[169]
                    }),
            .out_data(lut_168_out)
        );

reg   lut_168_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_168_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_168_ff <= lut_168_out;
    end
end

assign out_data[168] = lut_168_ff;




// LUT : 169

wire lut_169_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000010101010010101001110000000000000001000000110011000000110),
            .DEVICE(DEVICE)
        )
    i_lut_169
        (
            .in_data({
                         in_data[237],
                         in_data[1010],
                         in_data[557],
                         in_data[782],
                         in_data[85],
                         in_data[761]
                    }),
            .out_data(lut_169_out)
        );

reg   lut_169_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_169_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_169_ff <= lut_169_out;
    end
end

assign out_data[169] = lut_169_ff;




// LUT : 170

wire lut_170_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101110101010111111110111101111101111001110111111111100110011),
            .DEVICE(DEVICE)
        )
    i_lut_170
        (
            .in_data({
                         in_data[803],
                         in_data[894],
                         in_data[404],
                         in_data[388],
                         in_data[833],
                         in_data[543]
                    }),
            .out_data(lut_170_out)
        );

reg   lut_170_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_170_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_170_ff <= lut_170_out;
    end
end

assign out_data[170] = lut_170_ff;




// LUT : 171

wire lut_171_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000000000010011101011001000100000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_171
        (
            .in_data({
                         in_data[290],
                         in_data[57],
                         in_data[55],
                         in_data[798],
                         in_data[565],
                         in_data[21]
                    }),
            .out_data(lut_171_out)
        );

reg   lut_171_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_171_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_171_ff <= lut_171_out;
    end
end

assign out_data[171] = lut_171_ff;




// LUT : 172

wire lut_172_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000000100101010000000100000001110000011000000),
            .DEVICE(DEVICE)
        )
    i_lut_172
        (
            .in_data({
                         in_data[722],
                         in_data[683],
                         in_data[1005],
                         in_data[1018],
                         in_data[79],
                         in_data[799]
                    }),
            .out_data(lut_172_out)
        );

reg   lut_172_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_172_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_172_ff <= lut_172_out;
    end
end

assign out_data[172] = lut_172_ff;




// LUT : 173

wire lut_173_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100000010000000110000000000011111011010100010001000000010000),
            .DEVICE(DEVICE)
        )
    i_lut_173
        (
            .in_data({
                         in_data[422],
                         in_data[31],
                         in_data[145],
                         in_data[548],
                         in_data[546],
                         in_data[555]
                    }),
            .out_data(lut_173_out)
        );

reg   lut_173_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_173_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_173_ff <= lut_173_out;
    end
end

assign out_data[173] = lut_173_ff;




// LUT : 174

wire lut_174_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101000000010100100110000000100001010000100100000110100010000),
            .DEVICE(DEVICE)
        )
    i_lut_174
        (
            .in_data({
                         in_data[897],
                         in_data[243],
                         in_data[765],
                         in_data[185],
                         in_data[296],
                         in_data[380]
                    }),
            .out_data(lut_174_out)
        );

reg   lut_174_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_174_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_174_ff <= lut_174_out;
    end
end

assign out_data[174] = lut_174_ff;




// LUT : 175

wire lut_175_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111011111111111111111111111111011000111110101100100011111010),
            .DEVICE(DEVICE)
        )
    i_lut_175
        (
            .in_data({
                         in_data[341],
                         in_data[67],
                         in_data[38],
                         in_data[830],
                         in_data[532],
                         in_data[1017]
                    }),
            .out_data(lut_175_out)
        );

reg   lut_175_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_175_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_175_ff <= lut_175_out;
    end
end

assign out_data[175] = lut_175_ff;




// LUT : 176

wire lut_176_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110111110111111111111111111111111111111111111111111010111110100),
            .DEVICE(DEVICE)
        )
    i_lut_176
        (
            .in_data({
                         in_data[431],
                         in_data[349],
                         in_data[590],
                         in_data[343],
                         in_data[392],
                         in_data[427]
                    }),
            .out_data(lut_176_out)
        );

reg   lut_176_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_176_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_176_ff <= lut_176_out;
    end
end

assign out_data[176] = lut_176_ff;




// LUT : 177

wire lut_177_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110000000000111001110111010100010001000000010111010001110100),
            .DEVICE(DEVICE)
        )
    i_lut_177
        (
            .in_data({
                         in_data[701],
                         in_data[716],
                         in_data[391],
                         in_data[920],
                         in_data[698],
                         in_data[76]
                    }),
            .out_data(lut_177_out)
        );

reg   lut_177_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_177_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_177_ff <= lut_177_out;
    end
end

assign out_data[177] = lut_177_ff;




// LUT : 178

wire lut_178_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111011111111111111101111110001110100011111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_178
        (
            .in_data({
                         in_data[133],
                         in_data[294],
                         in_data[593],
                         in_data[682],
                         in_data[110],
                         in_data[466]
                    }),
            .out_data(lut_178_out)
        );

reg   lut_178_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_178_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_178_ff <= lut_178_out;
    end
end

assign out_data[178] = lut_178_ff;




// LUT : 179

wire lut_179_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011101011101100111010001110111111011111111111111111101011111),
            .DEVICE(DEVICE)
        )
    i_lut_179
        (
            .in_data({
                         in_data[695],
                         in_data[10],
                         in_data[553],
                         in_data[409],
                         in_data[436],
                         in_data[530]
                    }),
            .out_data(lut_179_out)
        );

reg   lut_179_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_179_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_179_ff <= lut_179_out;
    end
end

assign out_data[179] = lut_179_ff;




// LUT : 180

wire lut_180_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110011001100001110000001000011111110111011100011111000000000),
            .DEVICE(DEVICE)
        )
    i_lut_180
        (
            .in_data({
                         in_data[868],
                         in_data[696],
                         in_data[623],
                         in_data[470],
                         in_data[579],
                         in_data[651]
                    }),
            .out_data(lut_180_out)
        );

reg   lut_180_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_180_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_180_ff <= lut_180_out;
    end
end

assign out_data[180] = lut_180_ff;




// LUT : 181

wire lut_181_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110000000000000000000000000010111000111100000000010101101001),
            .DEVICE(DEVICE)
        )
    i_lut_181
        (
            .in_data({
                         in_data[521],
                         in_data[788],
                         in_data[386],
                         in_data[199],
                         in_data[805],
                         in_data[554]
                    }),
            .out_data(lut_181_out)
        );

reg   lut_181_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_181_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_181_ff <= lut_181_out;
    end
end

assign out_data[181] = lut_181_ff;




// LUT : 182

wire lut_182_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110100010111111111110011111110101001000101111011111110111),
            .DEVICE(DEVICE)
        )
    i_lut_182
        (
            .in_data({
                         in_data[174],
                         in_data[148],
                         in_data[966],
                         in_data[729],
                         in_data[820],
                         in_data[755]
                    }),
            .out_data(lut_182_out)
        );

reg   lut_182_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_182_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_182_ff <= lut_182_out;
    end
end

assign out_data[182] = lut_182_ff;




// LUT : 183

wire lut_183_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111101111111010111111111111111111111111111110101111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_183
        (
            .in_data({
                         in_data[280],
                         in_data[904],
                         in_data[501],
                         in_data[285],
                         in_data[777],
                         in_data[717]
                    }),
            .out_data(lut_183_out)
        );

reg   lut_183_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_183_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_183_ff <= lut_183_out;
    end
end

assign out_data[183] = lut_183_ff;




// LUT : 184

wire lut_184_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111011100000111010101100000011111111111011111111110011000000),
            .DEVICE(DEVICE)
        )
    i_lut_184
        (
            .in_data({
                         in_data[747],
                         in_data[1001],
                         in_data[162],
                         in_data[314],
                         in_data[457],
                         in_data[410]
                    }),
            .out_data(lut_184_out)
        );

reg   lut_184_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_184_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_184_ff <= lut_184_out;
    end
end

assign out_data[184] = lut_184_ff;




// LUT : 185

wire lut_185_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001000110000110100001111000000110011101100010011000110110001),
            .DEVICE(DEVICE)
        )
    i_lut_185
        (
            .in_data({
                         in_data[315],
                         in_data[784],
                         in_data[525],
                         in_data[520],
                         in_data[943],
                         in_data[464]
                    }),
            .out_data(lut_185_out)
        );

reg   lut_185_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_185_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_185_ff <= lut_185_out;
    end
end

assign out_data[185] = lut_185_ff;




// LUT : 186

wire lut_186_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101010001000000110111010111101100101000000000111011111110001),
            .DEVICE(DEVICE)
        )
    i_lut_186
        (
            .in_data({
                         in_data[146],
                         in_data[22],
                         in_data[104],
                         in_data[577],
                         in_data[331],
                         in_data[500]
                    }),
            .out_data(lut_186_out)
        );

reg   lut_186_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_186_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_186_ff <= lut_186_out;
    end
end

assign out_data[186] = lut_186_ff;




// LUT : 187

wire lut_187_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011101100000101101000100000000010111010010111110000001000000010),
            .DEVICE(DEVICE)
        )
    i_lut_187
        (
            .in_data({
                         in_data[203],
                         in_data[108],
                         in_data[774],
                         in_data[689],
                         in_data[488],
                         in_data[571]
                    }),
            .out_data(lut_187_out)
        );

reg   lut_187_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_187_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_187_ff <= lut_187_out;
    end
end

assign out_data[187] = lut_187_ff;




// LUT : 188

wire lut_188_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001111111111001110111011111100000100000001100110001111000111),
            .DEVICE(DEVICE)
        )
    i_lut_188
        (
            .in_data({
                         in_data[212],
                         in_data[712],
                         in_data[738],
                         in_data[169],
                         in_data[923],
                         in_data[113]
                    }),
            .out_data(lut_188_out)
        );

reg   lut_188_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_188_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_188_ff <= lut_188_out;
    end
end

assign out_data[188] = lut_188_ff;




// LUT : 189

wire lut_189_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101100001000000111000000110011101111000000001110110010000100),
            .DEVICE(DEVICE)
        )
    i_lut_189
        (
            .in_data({
                         in_data[5],
                         in_data[710],
                         in_data[821],
                         in_data[44],
                         in_data[676],
                         in_data[970]
                    }),
            .out_data(lut_189_out)
        );

reg   lut_189_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_189_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_189_ff <= lut_189_out;
    end
end

assign out_data[189] = lut_189_ff;




// LUT : 190

wire lut_190_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100001100000110000001100000011001110111011001100100011001000),
            .DEVICE(DEVICE)
        )
    i_lut_190
        (
            .in_data({
                         in_data[428],
                         in_data[196],
                         in_data[230],
                         in_data[604],
                         in_data[601],
                         in_data[924]
                    }),
            .out_data(lut_190_out)
        );

reg   lut_190_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_190_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_190_ff <= lut_190_out;
    end
end

assign out_data[190] = lut_190_ff;




// LUT : 191

wire lut_191_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110111111111111111111111100001100111011101100110111111111),
            .DEVICE(DEVICE)
        )
    i_lut_191
        (
            .in_data({
                         in_data[398],
                         in_data[127],
                         in_data[592],
                         in_data[862],
                         in_data[935],
                         in_data[890]
                    }),
            .out_data(lut_191_out)
        );

reg   lut_191_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_191_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_191_ff <= lut_191_out;
    end
end

assign out_data[191] = lut_191_ff;




// LUT : 192

wire lut_192_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000100000000000000010000000000000000000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_192
        (
            .in_data({
                         in_data[569],
                         in_data[68],
                         in_data[403],
                         in_data[492],
                         in_data[824],
                         in_data[235]
                    }),
            .out_data(lut_192_out)
        );

reg   lut_192_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_192_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_192_ff <= lut_192_out;
    end
end

assign out_data[192] = lut_192_ff;




// LUT : 193

wire lut_193_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000110010001111100011101000111111101111111111110010001100110011),
            .DEVICE(DEVICE)
        )
    i_lut_193
        (
            .in_data({
                         in_data[754],
                         in_data[641],
                         in_data[423],
                         in_data[936],
                         in_data[535],
                         in_data[111]
                    }),
            .out_data(lut_193_out)
        );

reg   lut_193_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_193_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_193_ff <= lut_193_out;
    end
end

assign out_data[193] = lut_193_ff;




// LUT : 194

wire lut_194_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111111111111110101010101111111010111111111110101010100000101),
            .DEVICE(DEVICE)
        )
    i_lut_194
        (
            .in_data({
                         in_data[390],
                         in_data[782],
                         in_data[853],
                         in_data[587],
                         in_data[572],
                         in_data[107]
                    }),
            .out_data(lut_194_out)
        );

reg   lut_194_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_194_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_194_ff <= lut_194_out;
    end
end

assign out_data[194] = lut_194_ff;




// LUT : 195

wire lut_195_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011101010110010100000000000000010111010101111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_195
        (
            .in_data({
                         in_data[887],
                         in_data[159],
                         in_data[510],
                         in_data[81],
                         in_data[4],
                         in_data[997]
                    }),
            .out_data(lut_195_out)
        );

reg   lut_195_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_195_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_195_ff <= lut_195_out;
    end
end

assign out_data[195] = lut_195_ff;




// LUT : 196

wire lut_196_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000001010101000000000010000011110001110100010111000100010000),
            .DEVICE(DEVICE)
        )
    i_lut_196
        (
            .in_data({
                         in_data[304],
                         in_data[255],
                         in_data[522],
                         in_data[401],
                         in_data[829],
                         in_data[780]
                    }),
            .out_data(lut_196_out)
        );

reg   lut_196_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_196_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_196_ff <= lut_196_out;
    end
end

assign out_data[196] = lut_196_ff;




// LUT : 197

wire lut_197_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000011111101110011111111111111001101111111111111111101111111),
            .DEVICE(DEVICE)
        )
    i_lut_197
        (
            .in_data({
                         in_data[1004],
                         in_data[700],
                         in_data[480],
                         in_data[463],
                         in_data[298],
                         in_data[197]
                    }),
            .out_data(lut_197_out)
        );

reg   lut_197_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_197_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_197_ff <= lut_197_out;
    end
end

assign out_data[197] = lut_197_ff;




// LUT : 198

wire lut_198_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000000010001000000000001000101000000000100010001000010010001),
            .DEVICE(DEVICE)
        )
    i_lut_198
        (
            .in_data({
                         in_data[96],
                         in_data[711],
                         in_data[783],
                         in_data[737],
                         in_data[511],
                         in_data[178]
                    }),
            .out_data(lut_198_out)
        );

reg   lut_198_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_198_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_198_ff <= lut_198_out;
    end
end

assign out_data[198] = lut_198_ff;




// LUT : 199

wire lut_199_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111110111111100111111001111111111111111111111001111111111),
            .DEVICE(DEVICE)
        )
    i_lut_199
        (
            .in_data({
                         in_data[541],
                         in_data[552],
                         in_data[418],
                         in_data[35],
                         in_data[26],
                         in_data[1009]
                    }),
            .out_data(lut_199_out)
        );

reg   lut_199_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_199_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_199_ff <= lut_199_out;
    end
end

assign out_data[199] = lut_199_ff;




// LUT : 200

wire lut_200_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000010110011000100010001011100000110111110111101000000),
            .DEVICE(DEVICE)
        )
    i_lut_200
        (
            .in_data({
                         in_data[503],
                         in_data[596],
                         in_data[969],
                         in_data[92],
                         in_data[97],
                         in_data[496]
                    }),
            .out_data(lut_200_out)
        );

reg   lut_200_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_200_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_200_ff <= lut_200_out;
    end
end

assign out_data[200] = lut_200_ff;




// LUT : 201

wire lut_201_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001111110010010100111111101111110000111110111110111111111010),
            .DEVICE(DEVICE)
        )
    i_lut_201
        (
            .in_data({
                         in_data[670],
                         in_data[381],
                         in_data[49],
                         in_data[58],
                         in_data[815],
                         in_data[907]
                    }),
            .out_data(lut_201_out)
        );

reg   lut_201_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_201_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_201_ff <= lut_201_out;
    end
end

assign out_data[201] = lut_201_ff;




// LUT : 202

wire lut_202_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010100001101000000000100000000000000010100000101101000001111000),
            .DEVICE(DEVICE)
        )
    i_lut_202
        (
            .in_data({
                         in_data[507],
                         in_data[516],
                         in_data[177],
                         in_data[346],
                         in_data[804],
                         in_data[369]
                    }),
            .out_data(lut_202_out)
        );

reg   lut_202_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_202_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_202_ff <= lut_202_out;
    end
end

assign out_data[202] = lut_202_ff;




// LUT : 203

wire lut_203_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010100011110010010000100110100100010111111100100010101011111),
            .DEVICE(DEVICE)
        )
    i_lut_203
        (
            .in_data({
                         in_data[80],
                         in_data[53],
                         in_data[479],
                         in_data[878],
                         in_data[359],
                         in_data[678]
                    }),
            .out_data(lut_203_out)
        );

reg   lut_203_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_203_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_203_ff <= lut_203_out;
    end
end

assign out_data[203] = lut_203_ff;




// LUT : 204

wire lut_204_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100010011110111000000001010000011110100111101111101000011100100),
            .DEVICE(DEVICE)
        )
    i_lut_204
        (
            .in_data({
                         in_data[929],
                         in_data[261],
                         in_data[752],
                         in_data[908],
                         in_data[812],
                         in_data[732]
                    }),
            .out_data(lut_204_out)
        );

reg   lut_204_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_204_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_204_ff <= lut_204_out;
    end
end

assign out_data[204] = lut_204_ff;




// LUT : 205

wire lut_205_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001111111111111111111111111111011111111111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_205
        (
            .in_data({
                         in_data[808],
                         in_data[508],
                         in_data[94],
                         in_data[705],
                         in_data[807],
                         in_data[687]
                    }),
            .out_data(lut_205_out)
        );

reg   lut_205_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_205_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_205_ff <= lut_205_out;
    end
end

assign out_data[205] = lut_205_ff;




// LUT : 206

wire lut_206_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001111111111111101111111111111111111111111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_206
        (
            .in_data({
                         in_data[588],
                         in_data[991],
                         in_data[911],
                         in_data[143],
                         in_data[512],
                         in_data[615]
                    }),
            .out_data(lut_206_out)
        );

reg   lut_206_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_206_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_206_ff <= lut_206_out;
    end
end

assign out_data[206] = lut_206_ff;




// LUT : 207

wire lut_207_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010111011111000000010101110100000000011111110001000001010101),
            .DEVICE(DEVICE)
        )
    i_lut_207
        (
            .in_data({
                         in_data[677],
                         in_data[414],
                         in_data[364],
                         in_data[801],
                         in_data[240],
                         in_data[865]
                    }),
            .out_data(lut_207_out)
        );

reg   lut_207_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_207_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_207_ff <= lut_207_out;
    end
end

assign out_data[207] = lut_207_ff;




// LUT : 208

wire lut_208_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110000010000000111110000000001001100000000000100110101000100),
            .DEVICE(DEVICE)
        )
    i_lut_208
        (
            .in_data({
                         in_data[291],
                         in_data[665],
                         in_data[362],
                         in_data[888],
                         in_data[472],
                         in_data[919]
                    }),
            .out_data(lut_208_out)
        );

reg   lut_208_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_208_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_208_ff <= lut_208_out;
    end
end

assign out_data[208] = lut_208_ff;




// LUT : 209

wire lut_209_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101111101100111110111100100011111111111011001111111111001100),
            .DEVICE(DEVICE)
        )
    i_lut_209
        (
            .in_data({
                         in_data[241],
                         in_data[217],
                         in_data[487],
                         in_data[282],
                         in_data[312],
                         in_data[206]
                    }),
            .out_data(lut_209_out)
        );

reg   lut_209_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_209_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_209_ff <= lut_209_out;
    end
end

assign out_data[209] = lut_209_ff;




// LUT : 210

wire lut_210_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000001000000000000010001110111100000000010001100),
            .DEVICE(DEVICE)
        )
    i_lut_210
        (
            .in_data({
                         in_data[112],
                         in_data[947],
                         in_data[211],
                         in_data[713],
                         in_data[618],
                         in_data[645]
                    }),
            .out_data(lut_210_out)
        );

reg   lut_210_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_210_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_210_ff <= lut_210_out;
    end
end

assign out_data[210] = lut_210_ff;




// LUT : 211

wire lut_211_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111110111010101001011110001110111011101010000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_211
        (
            .in_data({
                         in_data[417],
                         in_data[297],
                         in_data[256],
                         in_data[895],
                         in_data[855],
                         in_data[134]
                    }),
            .out_data(lut_211_out)
        );

reg   lut_211_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_211_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_211_ff <= lut_211_out;
    end
end

assign out_data[211] = lut_211_ff;




// LUT : 212

wire lut_212_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000011101111101111001111111101111111111111111111111110111111),
            .DEVICE(DEVICE)
        )
    i_lut_212
        (
            .in_data({
                         in_data[485],
                         in_data[836],
                         in_data[330],
                         in_data[674],
                         in_data[956],
                         in_data[220]
                    }),
            .out_data(lut_212_out)
        );

reg   lut_212_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_212_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_212_ff <= lut_212_out;
    end
end

assign out_data[212] = lut_212_ff;




// LUT : 213

wire lut_213_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100100000001010100000000000101000001000000010000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_213
        (
            .in_data({
                         in_data[41],
                         in_data[961],
                         in_data[168],
                         in_data[411],
                         in_data[514],
                         in_data[809]
                    }),
            .out_data(lut_213_out)
        );

reg   lut_213_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_213_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_213_ff <= lut_213_out;
    end
end

assign out_data[213] = lut_213_ff;




// LUT : 214

wire lut_214_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111011111111111000001011111111110110000110001011111100010110010),
            .DEVICE(DEVICE)
        )
    i_lut_214
        (
            .in_data({
                         in_data[896],
                         in_data[575],
                         in_data[126],
                         in_data[558],
                         in_data[599],
                         in_data[685]
                    }),
            .out_data(lut_214_out)
        );

reg   lut_214_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_214_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_214_ff <= lut_214_out;
    end
end

assign out_data[214] = lut_214_ff;




// LUT : 215

wire lut_215_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101110000111010111110101111111011101000000001111111100010011),
            .DEVICE(DEVICE)
        )
    i_lut_215
        (
            .in_data({
                         in_data[356],
                         in_data[556],
                         in_data[263],
                         in_data[257],
                         in_data[19],
                         in_data[629]
                    }),
            .out_data(lut_215_out)
        );

reg   lut_215_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_215_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_215_ff <= lut_215_out;
    end
end

assign out_data[215] = lut_215_ff;




// LUT : 216

wire lut_216_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010100000000111111110000000011010100001000001111111100000000),
            .DEVICE(DEVICE)
        )
    i_lut_216
        (
            .in_data({
                         in_data[320],
                         in_data[594],
                         in_data[59],
                         in_data[946],
                         in_data[46],
                         in_data[994]
                    }),
            .out_data(lut_216_out)
        );

reg   lut_216_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_216_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_216_ff <= lut_216_out;
    end
end

assign out_data[216] = lut_216_ff;




// LUT : 217

wire lut_217_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000111010101010100011101011101000000000000001101000011010100),
            .DEVICE(DEVICE)
        )
    i_lut_217
        (
            .in_data({
                         in_data[15],
                         in_data[714],
                         in_data[375],
                         in_data[1021],
                         in_data[276],
                         in_data[750]
                    }),
            .out_data(lut_217_out)
        );

reg   lut_217_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_217_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_217_ff <= lut_217_out;
    end
end

assign out_data[217] = lut_217_ff;




// LUT : 218

wire lut_218_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010100000000011101111001000000000101000000001101110101100101),
            .DEVICE(DEVICE)
        )
    i_lut_218
        (
            .in_data({
                         in_data[948],
                         in_data[998],
                         in_data[574],
                         in_data[1006],
                         in_data[336],
                         in_data[976]
                    }),
            .out_data(lut_218_out)
        );

reg   lut_218_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_218_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_218_ff <= lut_218_out;
    end
end

assign out_data[218] = lut_218_ff;




// LUT : 219

wire lut_219_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111011111111111111101111011111111110111011111111011011000),
            .DEVICE(DEVICE)
        )
    i_lut_219
        (
            .in_data({
                         in_data[218],
                         in_data[529],
                         in_data[1016],
                         in_data[308],
                         in_data[65],
                         in_data[658]
                    }),
            .out_data(lut_219_out)
        );

reg   lut_219_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_219_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_219_ff <= lut_219_out;
    end
end

assign out_data[219] = lut_219_ff;




// LUT : 220

wire lut_220_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101011000000101110101110101000000000010000000000100001000000),
            .DEVICE(DEVICE)
        )
    i_lut_220
        (
            .in_data({
                         in_data[958],
                         in_data[668],
                         in_data[892],
                         in_data[254],
                         in_data[78],
                         in_data[771]
                    }),
            .out_data(lut_220_out)
        );

reg   lut_220_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_220_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_220_ff <= lut_220_out;
    end
end

assign out_data[220] = lut_220_ff;




// LUT : 221

wire lut_221_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000000100000000000000000001011101010111011001100000011000000),
            .DEVICE(DEVICE)
        )
    i_lut_221
        (
            .in_data({
                         in_data[724],
                         in_data[29],
                         in_data[216],
                         in_data[775],
                         in_data[426],
                         in_data[497]
                    }),
            .out_data(lut_221_out)
        );

reg   lut_221_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_221_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_221_ff <= lut_221_out;
    end
end

assign out_data[221] = lut_221_ff;




// LUT : 222

wire lut_222_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000000000000010100100010111101110001000000000111011101110111),
            .DEVICE(DEVICE)
        )
    i_lut_222
        (
            .in_data({
                         in_data[232],
                         in_data[719],
                         in_data[609],
                         in_data[299],
                         in_data[453],
                         in_data[768]
                    }),
            .out_data(lut_222_out)
        );

reg   lut_222_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_222_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_222_ff <= lut_222_out;
    end
end

assign out_data[222] = lut_222_ff;




// LUT : 223

wire lut_223_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001100100010111111110011001100110111000101110111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_223
        (
            .in_data({
                         in_data[225],
                         in_data[277],
                         in_data[286],
                         in_data[440],
                         in_data[916],
                         in_data[886]
                    }),
            .out_data(lut_223_out)
        );

reg   lut_223_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_223_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_223_ff <= lut_223_out;
    end
end

assign out_data[223] = lut_223_ff;




// LUT : 224

wire lut_224_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111100110011000000110000001100110101000001010000001100000001),
            .DEVICE(DEVICE)
        )
    i_lut_224
        (
            .in_data({
                         in_data[989],
                         in_data[980],
                         in_data[325],
                         in_data[523],
                         in_data[628],
                         in_data[419]
                    }),
            .out_data(lut_224_out)
        );

reg   lut_224_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_224_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_224_ff <= lut_224_out;
    end
end

assign out_data[224] = lut_224_ff;




// LUT : 225

wire lut_225_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000111110101111111011111111100010100011101010101011100110000),
            .DEVICE(DEVICE)
        )
    i_lut_225
        (
            .in_data({
                         in_data[746],
                         in_data[33],
                         in_data[438],
                         in_data[983],
                         in_data[1000],
                         in_data[1019]
                    }),
            .out_data(lut_225_out)
        );

reg   lut_225_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_225_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_225_ff <= lut_225_out;
    end
end

assign out_data[225] = lut_225_ff;




// LUT : 226

wire lut_226_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101000001010000000001011011100101010101110011010011011111100),
            .DEVICE(DEVICE)
        )
    i_lut_226
        (
            .in_data({
                         in_data[355],
                         in_data[478],
                         in_data[114],
                         in_data[933],
                         in_data[115],
                         in_data[242]
                    }),
            .out_data(lut_226_out)
        );

reg   lut_226_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_226_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_226_ff <= lut_226_out;
    end
end

assign out_data[226] = lut_226_ff;




// LUT : 227

wire lut_227_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110111111100110111011011101011111111111100000111111111000000),
            .DEVICE(DEVICE)
        )
    i_lut_227
        (
            .in_data({
                         in_data[509],
                         in_data[938],
                         in_data[876],
                         in_data[723],
                         in_data[213],
                         in_data[733]
                    }),
            .out_data(lut_227_out)
        );

reg   lut_227_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_227_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_227_ff <= lut_227_out;
    end
end

assign out_data[227] = lut_227_ff;




// LUT : 228

wire lut_228_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101001001010000011010110000000001100010010100000011001100110010),
            .DEVICE(DEVICE)
        )
    i_lut_228
        (
            .in_data({
                         in_data[1014],
                         in_data[550],
                         in_data[47],
                         in_data[400],
                         in_data[643],
                         in_data[880]
                    }),
            .out_data(lut_228_out)
        );

reg   lut_228_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_228_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_228_ff <= lut_228_out;
    end
end

assign out_data[228] = lut_228_ff;




// LUT : 229

wire lut_229_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111110111111001011110010111111111111111111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_229
        (
            .in_data({
                         in_data[365],
                         in_data[531],
                         in_data[597],
                         in_data[840],
                         in_data[959],
                         in_data[627]
                    }),
            .out_data(lut_229_out)
        );

reg   lut_229_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_229_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_229_ff <= lut_229_out;
    end
end

assign out_data[229] = lut_229_ff;




// LUT : 230

wire lut_230_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101011000110011110111001011101010000000000000101000100010101),
            .DEVICE(DEVICE)
        )
    i_lut_230
        (
            .in_data({
                         in_data[679],
                         in_data[591],
                         in_data[222],
                         in_data[20],
                         in_data[690],
                         in_data[1020]
                    }),
            .out_data(lut_230_out)
        );

reg   lut_230_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_230_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_230_ff <= lut_230_out;
    end
end

assign out_data[230] = lut_230_ff;




// LUT : 231

wire lut_231_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000000000000010100010000000000000000000000010),
            .DEVICE(DEVICE)
        )
    i_lut_231
        (
            .in_data({
                         in_data[666],
                         in_data[189],
                         in_data[382],
                         in_data[173],
                         in_data[759],
                         in_data[505]
                    }),
            .out_data(lut_231_out)
        );

reg   lut_231_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_231_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_231_ff <= lut_231_out;
    end
end

assign out_data[231] = lut_231_ff;




// LUT : 232

wire lut_232_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010100001101000000000000100000000100000001000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_232
        (
            .in_data({
                         in_data[495],
                         in_data[156],
                         in_data[963],
                         in_data[644],
                         in_data[937],
                         in_data[132]
                    }),
            .out_data(lut_232_out)
        );

reg   lut_232_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_232_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_232_ff <= lut_232_out;
    end
end

assign out_data[232] = lut_232_ff;




// LUT : 233

wire lut_233_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000110000000101000010011010000000000000000100001000000000),
            .DEVICE(DEVICE)
        )
    i_lut_233
        (
            .in_data({
                         in_data[373],
                         in_data[367],
                         in_data[939],
                         in_data[128],
                         in_data[684],
                         in_data[284]
                    }),
            .out_data(lut_233_out)
        );

reg   lut_233_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_233_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_233_ff <= lut_233_out;
    end
end

assign out_data[233] = lut_233_ff;




// LUT : 234

wire lut_234_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111100111111011111110011111111111101111111101111111011111111),
            .DEVICE(DEVICE)
        )
    i_lut_234
        (
            .in_data({
                         in_data[761],
                         in_data[141],
                         in_data[625],
                         in_data[361],
                         in_data[631],
                         in_data[582]
                    }),
            .out_data(lut_234_out)
        );

reg   lut_234_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_234_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_234_ff <= lut_234_out;
    end
end

assign out_data[234] = lut_234_ff;




// LUT : 235

wire lut_235_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000011110000111100111111001111111011111100011111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_235
        (
            .in_data({
                         in_data[194],
                         in_data[871],
                         in_data[420],
                         in_data[433],
                         in_data[832],
                         in_data[730]
                    }),
            .out_data(lut_235_out)
        );

reg   lut_235_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_235_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_235_ff <= lut_235_out;
    end
end

assign out_data[235] = lut_235_ff;




// LUT : 236

wire lut_236_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101110101111101011111011110110000011011011011111100110111001100),
            .DEVICE(DEVICE)
        )
    i_lut_236
        (
            .in_data({
                         in_data[718],
                         in_data[233],
                         in_data[62],
                         in_data[321],
                         in_data[71],
                         in_data[973]
                    }),
            .out_data(lut_236_out)
        );

reg   lut_236_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_236_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_236_ff <= lut_236_out;
    end
end

assign out_data[236] = lut_236_ff;




// LUT : 237

wire lut_237_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110100001000111001001111011000010101000001010000000000100000),
            .DEVICE(DEVICE)
        )
    i_lut_237
        (
            .in_data({
                         in_data[639],
                         in_data[726],
                         in_data[316],
                         in_data[376],
                         in_data[228],
                         in_data[751]
                    }),
            .out_data(lut_237_out)
        );

reg   lut_237_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_237_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_237_ff <= lut_237_out;
    end
end

assign out_data[237] = lut_237_ff;




// LUT : 238

wire lut_238_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110101110111111111111111111111111111011101111111111111100),
            .DEVICE(DEVICE)
        )
    i_lut_238
        (
            .in_data({
                         in_data[374],
                         in_data[842],
                         in_data[90],
                         in_data[773],
                         in_data[252],
                         in_data[142]
                    }),
            .out_data(lut_238_out)
        );

reg   lut_238_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_238_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_238_ff <= lut_238_out;
    end
end

assign out_data[238] = lut_238_ff;




// LUT : 239

wire lut_239_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001000000000000001101000000000010010010000000001011001100),
            .DEVICE(DEVICE)
        )
    i_lut_239
        (
            .in_data({
                         in_data[278],
                         in_data[75],
                         in_data[48],
                         in_data[292],
                         in_data[180],
                         in_data[149]
                    }),
            .out_data(lut_239_out)
        );

reg   lut_239_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_239_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_239_ff <= lut_239_out;
    end
end

assign out_data[239] = lut_239_ff;




// LUT : 240

wire lut_240_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110011111100111111011111110100111100010101000001000101010101),
            .DEVICE(DEVICE)
        )
    i_lut_240
        (
            .in_data({
                         in_data[397],
                         in_data[125],
                         in_data[536],
                         in_data[952],
                         in_data[279],
                         in_data[319]
                    }),
            .out_data(lut_240_out)
        );

reg   lut_240_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_240_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_240_ff <= lut_240_out;
    end
end

assign out_data[240] = lut_240_ff;




// LUT : 241

wire lut_241_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111101110011000000110000000000110011001100110000001100000010),
            .DEVICE(DEVICE)
        )
    i_lut_241
        (
            .in_data({
                         in_data[221],
                         in_data[881],
                         in_data[557],
                         in_data[638],
                         in_data[694],
                         in_data[534]
                    }),
            .out_data(lut_241_out)
        );

reg   lut_241_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_241_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_241_ff <= lut_241_out;
    end
end

assign out_data[241] = lut_241_ff;




// LUT : 242

wire lut_242_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000001110000011111111111100000000000010100010011111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_242
        (
            .in_data({
                         in_data[838],
                         in_data[883],
                         in_data[253],
                         in_data[482],
                         in_data[987],
                         in_data[144]
                    }),
            .out_data(lut_242_out)
        );

reg   lut_242_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_242_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_242_ff <= lut_242_out;
    end
end

assign out_data[242] = lut_242_ff;




// LUT : 243

wire lut_243_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111100000000000001000000000010110000000000010000000000000011),
            .DEVICE(DEVICE)
        )
    i_lut_243
        (
            .in_data({
                         in_data[105],
                         in_data[121],
                         in_data[318],
                         in_data[727],
                         in_data[721],
                         in_data[136]
                    }),
            .out_data(lut_243_out)
        );

reg   lut_243_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_243_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_243_ff <= lut_243_out;
    end
end

assign out_data[243] = lut_243_ff;




// LUT : 244

wire lut_244_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000010000010100000101010001000000000000001101000011111100),
            .DEVICE(DEVICE)
        )
    i_lut_244
        (
            .in_data({
                         in_data[826],
                         in_data[204],
                         in_data[657],
                         in_data[818],
                         in_data[456],
                         in_data[851]
                    }),
            .out_data(lut_244_out)
        );

reg   lut_244_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_244_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_244_ff <= lut_244_out;
    end
end

assign out_data[244] = lut_244_ff;




// LUT : 245

wire lut_245_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000110011110011010010101110001000000001100001000000000110100100),
            .DEVICE(DEVICE)
        )
    i_lut_245
        (
            .in_data({
                         in_data[934],
                         in_data[847],
                         in_data[300],
                         in_data[1010],
                         in_data[533],
                         in_data[849]
                    }),
            .out_data(lut_245_out)
        );

reg   lut_245_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_245_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_245_ff <= lut_245_out;
    end
end

assign out_data[245] = lut_245_ff;




// LUT : 246

wire lut_246_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000111100001010000111110101011000001100000011001110111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_246
        (
            .in_data({
                         in_data[25],
                         in_data[458],
                         in_data[675],
                         in_data[612],
                         in_data[673],
                         in_data[307]
                    }),
            .out_data(lut_246_out)
        );

reg   lut_246_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_246_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_246_ff <= lut_246_out;
    end
end

assign out_data[246] = lut_246_ff;




// LUT : 247

wire lut_247_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111101011011110111110101101100001101010011011100111100001101),
            .DEVICE(DEVICE)
        )
    i_lut_247
        (
            .in_data({
                         in_data[626],
                         in_data[633],
                         in_data[1015],
                         in_data[743],
                         in_data[607],
                         in_data[273]
                    }),
            .out_data(lut_247_out)
        );

reg   lut_247_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_247_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_247_ff <= lut_247_out;
    end
end

assign out_data[247] = lut_247_ff;




// LUT : 248

wire lut_248_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001001101000000000000000001000100010011010000100011000000110001),
            .DEVICE(DEVICE)
        )
    i_lut_248
        (
            .in_data({
                         in_data[342],
                         in_data[3],
                         in_data[14],
                         in_data[454],
                         in_data[451],
                         in_data[219]
                    }),
            .out_data(lut_248_out)
        );

reg   lut_248_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_248_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_248_ff <= lut_248_out;
    end
end

assign out_data[248] = lut_248_ff;




// LUT : 249

wire lut_249_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000000000000001000100000010000100010010100001010001001000100),
            .DEVICE(DEVICE)
        )
    i_lut_249
        (
            .in_data({
                         in_data[372],
                         in_data[899],
                         in_data[528],
                         in_data[210],
                         in_data[309],
                         in_data[234]
                    }),
            .out_data(lut_249_out)
        );

reg   lut_249_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_249_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_249_ff <= lut_249_out;
    end
end

assign out_data[249] = lut_249_ff;




// LUT : 250

wire lut_250_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010111111111110111011111110111110111111111011111110111011101),
            .DEVICE(DEVICE)
        )
    i_lut_250
        (
            .in_data({
                         in_data[161],
                         in_data[749],
                         in_data[944],
                         in_data[568],
                         in_data[745],
                         in_data[421]
                    }),
            .out_data(lut_250_out)
        );

reg   lut_250_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_250_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_250_ff <= lut_250_out;
    end
end

assign out_data[250] = lut_250_ff;




// LUT : 251

wire lut_251_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111101111111111111110100111010111111101110111110111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_251
        (
            .in_data({
                         in_data[953],
                         in_data[118],
                         in_data[82],
                         in_data[622],
                         in_data[340],
                         in_data[791]
                    }),
            .out_data(lut_251_out)
        );

reg   lut_251_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_251_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_251_ff <= lut_251_out;
    end
end

assign out_data[251] = lut_251_ff;




// LUT : 252

wire lut_252_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111111111111111111111111011100001001110111010101000111011101),
            .DEVICE(DEVICE)
        )
    i_lut_252
        (
            .in_data({
                         in_data[345],
                         in_data[659],
                         in_data[236],
                         in_data[461],
                         in_data[992],
                         in_data[109]
                    }),
            .out_data(lut_252_out)
        );

reg   lut_252_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_252_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_252_ff <= lut_252_out;
    end
end

assign out_data[252] = lut_252_ff;




// LUT : 253

wire lut_253_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011111011111110110101100100110011111111111111111111111111111100),
            .DEVICE(DEVICE)
        )
    i_lut_253
        (
            .in_data({
                         in_data[562],
                         in_data[123],
                         in_data[660],
                         in_data[184],
                         in_data[778],
                         in_data[301]
                    }),
            .out_data(lut_253_out)
        );

reg   lut_253_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_253_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_253_ff <= lut_253_out;
    end
end

assign out_data[253] = lut_253_ff;




// LUT : 254

wire lut_254_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000000000111001000000000001100100010001010110000000000000010),
            .DEVICE(DEVICE)
        )
    i_lut_254
        (
            .in_data({
                         in_data[407],
                         in_data[102],
                         in_data[692],
                         in_data[910],
                         in_data[990],
                         in_data[335]
                    }),
            .out_data(lut_254_out)
        );

reg   lut_254_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_254_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_254_ff <= lut_254_out;
    end
end

assign out_data[254] = lut_254_ff;




// LUT : 255

wire lut_255_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000100000000000000000000000000000100000000000000000010000000),
            .DEVICE(DEVICE)
        )
    i_lut_255
        (
            .in_data({
                         in_data[348],
                         in_data[786],
                         in_data[155],
                         in_data[439],
                         in_data[186],
                         in_data[691]
                    }),
            .out_data(lut_255_out)
        );

reg   lut_255_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_255_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_255_ff <= lut_255_out;
    end
end

assign out_data[255] = lut_255_ff;




// LUT : 256

wire lut_256_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1001010100011101111111011000100011111111111111101111110111111010),
            .DEVICE(DEVICE)
        )
    i_lut_256
        (
            .in_data({
                         in_data[954],
                         in_data[402],
                         in_data[905],
                         in_data[493],
                         in_data[515],
                         in_data[200]
                    }),
            .out_data(lut_256_out)
        );

reg   lut_256_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_256_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_256_ff <= lut_256_out;
    end
end

assign out_data[256] = lut_256_ff;




// LUT : 257

wire lut_257_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100111111011001010110010111111111101111101110010011100000101),
            .DEVICE(DEVICE)
        )
    i_lut_257
        (
            .in_data({
                         in_data[117],
                         in_data[408],
                         in_data[518],
                         in_data[913],
                         in_data[827],
                         in_data[352]
                    }),
            .out_data(lut_257_out)
        );

reg   lut_257_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_257_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_257_ff <= lut_257_out;
    end
end

assign out_data[257] = lut_257_ff;




// LUT : 258

wire lut_258_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001100101010010100111111111111100001000100000000010010100111110),
            .DEVICE(DEVICE)
        )
    i_lut_258
        (
            .in_data({
                         in_data[385],
                         in_data[1007],
                         in_data[964],
                         in_data[800],
                         in_data[739],
                         in_data[494]
                    }),
            .out_data(lut_258_out)
        );

reg   lut_258_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_258_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_258_ff <= lut_258_out;
    end
end

assign out_data[258] = lut_258_ff;




// LUT : 259

wire lut_259_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111111011101000001000000010000000000100010100000000000001100),
            .DEVICE(DEVICE)
        )
    i_lut_259
        (
            .in_data({
                         in_data[795],
                         in_data[925],
                         in_data[98],
                         in_data[150],
                         in_data[819],
                         in_data[450]
                    }),
            .out_data(lut_259_out)
        );

reg   lut_259_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_259_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_259_ff <= lut_259_out;
    end
end

assign out_data[259] = lut_259_ff;




// LUT : 260

wire lut_260_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000010100000111111000100000000000000000000001110100010000000),
            .DEVICE(DEVICE)
        )
    i_lut_260
        (
            .in_data({
                         in_data[559],
                         in_data[927],
                         in_data[789],
                         in_data[183],
                         in_data[560],
                         in_data[770]
                    }),
            .out_data(lut_260_out)
        );

reg   lut_260_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_260_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_260_ff <= lut_260_out;
    end
end

assign out_data[260] = lut_260_ff;




// LUT : 261

wire lut_261_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000100010000000000011101110100000001000100000001000110111),
            .DEVICE(DEVICE)
        )
    i_lut_261
        (
            .in_data({
                         in_data[51],
                         in_data[333],
                         in_data[227],
                         in_data[175],
                         in_data[37],
                         in_data[642]
                    }),
            .out_data(lut_261_out)
        );

reg   lut_261_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_261_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_261_ff <= lut_261_out;
    end
end

assign out_data[261] = lut_261_ff;




// LUT : 262

wire lut_262_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010100000000001101100000000001110001100011000111011010001000),
            .DEVICE(DEVICE)
        )
    i_lut_262
        (
            .in_data({
                         in_data[875],
                         in_data[858],
                         in_data[922],
                         in_data[247],
                         in_data[589],
                         in_data[311]
                    }),
            .out_data(lut_262_out)
        );

reg   lut_262_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_262_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_262_ff <= lut_262_out;
    end
end

assign out_data[262] = lut_262_ff;




// LUT : 263

wire lut_263_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111100000000111111111011001101011111101110111101111110111011),
            .DEVICE(DEVICE)
        )
    i_lut_263
        (
            .in_data({
                         in_data[167],
                         in_data[872],
                         in_data[606],
                         in_data[469],
                         in_data[583],
                         in_data[140]
                    }),
            .out_data(lut_263_out)
        );

reg   lut_263_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_263_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_263_ff <= lut_263_out;
    end
end

assign out_data[263] = lut_263_ff;




// LUT : 264

wire lut_264_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110111111111001100111110111111111111110011111010111000101110),
            .DEVICE(DEVICE)
        )
    i_lut_264
        (
            .in_data({
                         in_data[884],
                         in_data[1022],
                         in_data[416],
                         in_data[584],
                         in_data[776],
                         in_data[979]
                    }),
            .out_data(lut_264_out)
        );

reg   lut_264_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_264_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_264_ff <= lut_264_out;
    end
end

assign out_data[264] = lut_264_ff;




// LUT : 265

wire lut_265_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011111111111111111101110111111100010111101001110000011101100),
            .DEVICE(DEVICE)
        )
    i_lut_265
        (
            .in_data({
                         in_data[99],
                         in_data[813],
                         in_data[170],
                         in_data[347],
                         in_data[395],
                         in_data[344]
                    }),
            .out_data(lut_265_out)
        );

reg   lut_265_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_265_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_265_ff <= lut_265_out;
    end
end

assign out_data[265] = lut_265_ff;




// LUT : 266

wire lut_266_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101100000000000000100000001000000000000000000000000000001010),
            .DEVICE(DEVICE)
        )
    i_lut_266
        (
            .in_data({
                         in_data[915],
                         in_data[483],
                         in_data[8],
                         in_data[223],
                         in_data[708],
                         in_data[332]
                    }),
            .out_data(lut_266_out)
        );

reg   lut_266_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_266_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_266_ff <= lut_266_out;
    end
end

assign out_data[266] = lut_266_ff;




// LUT : 267

wire lut_267_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000001010101011011011100100011011000000001010111111101100),
            .DEVICE(DEVICE)
        )
    i_lut_267
        (
            .in_data({
                         in_data[368],
                         in_data[147],
                         in_data[655],
                         in_data[455],
                         in_data[753],
                         in_data[834]
                    }),
            .out_data(lut_267_out)
        );

reg   lut_267_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_267_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_267_ff <= lut_267_out;
    end
end

assign out_data[267] = lut_267_ff;




// LUT : 268

wire lut_268_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101000000000110000100000000000001111000001011100111100001101),
            .DEVICE(DEVICE)
        )
    i_lut_268
        (
            .in_data({
                         in_data[43],
                         in_data[36],
                         in_data[477],
                         in_data[328],
                         in_data[295],
                         in_data[860]
                    }),
            .out_data(lut_268_out)
        );

reg   lut_268_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_268_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_268_ff <= lut_268_out;
    end
end

assign out_data[268] = lut_268_ff;




// LUT : 269

wire lut_269_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000010000000110000101000000000000011010000001010101111),
            .DEVICE(DEVICE)
        )
    i_lut_269
        (
            .in_data({
                         in_data[163],
                         in_data[83],
                         in_data[846],
                         in_data[379],
                         in_data[837],
                         in_data[30]
                    }),
            .out_data(lut_269_out)
        );

reg   lut_269_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_269_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_269_ff <= lut_269_out;
    end
end

assign out_data[269] = lut_269_ff;




// LUT : 270

wire lut_270_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011110100010000001101010001000001011111000100110001110100010101),
            .DEVICE(DEVICE)
        )
    i_lut_270
        (
            .in_data({
                         in_data[506],
                         in_data[566],
                         in_data[215],
                         in_data[74],
                         in_data[322],
                         in_data[198]
                    }),
            .out_data(lut_270_out)
        );

reg   lut_270_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_270_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_270_ff <= lut_270_out;
    end
end

assign out_data[270] = lut_270_ff;




// LUT : 271

wire lut_271_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100000000100011000000000000001101000100001000000100010000000000),
            .DEVICE(DEVICE)
        )
    i_lut_271
        (
            .in_data({
                         in_data[467],
                         in_data[72],
                         in_data[489],
                         in_data[50],
                         in_data[731],
                         in_data[740]
                    }),
            .out_data(lut_271_out)
        );

reg   lut_271_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_271_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_271_ff <= lut_271_out;
    end
end

assign out_data[271] = lut_271_ff;




// LUT : 272

wire lut_272_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111101010000110000001000111011111100010000001010100010001000),
            .DEVICE(DEVICE)
        )
    i_lut_272
        (
            .in_data({
                         in_data[856],
                         in_data[757],
                         in_data[951],
                         in_data[524],
                         in_data[909],
                         in_data[993]
                    }),
            .out_data(lut_272_out)
        );

reg   lut_272_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_272_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_272_ff <= lut_272_out;
    end
end

assign out_data[272] = lut_272_ff;




// LUT : 273

wire lut_273_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111111111110111111111111101000011110000),
            .DEVICE(DEVICE)
        )
    i_lut_273
        (
            .in_data({
                         in_data[617],
                         in_data[100],
                         in_data[226],
                         in_data[984],
                         in_data[852],
                         in_data[637]
                    }),
            .out_data(lut_273_out)
        );

reg   lut_273_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_273_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_273_ff <= lut_273_out;
    end
end

assign out_data[273] = lut_273_ff;




// LUT : 274

wire lut_274_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001111111111010001001000000011110010111100001110110001100100),
            .DEVICE(DEVICE)
        )
    i_lut_274
        (
            .in_data({
                         in_data[706],
                         in_data[0],
                         in_data[867],
                         in_data[975],
                         in_data[527],
                         in_data[13]
                    }),
            .out_data(lut_274_out)
        );

reg   lut_274_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_274_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_274_ff <= lut_274_out;
    end
end

assign out_data[274] = lut_274_ff;




// LUT : 275

wire lut_275_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000000000000010000000000000011100111111011100110010010000010),
            .DEVICE(DEVICE)
        )
    i_lut_275
        (
            .in_data({
                         in_data[244],
                         in_data[828],
                         in_data[649],
                         in_data[12],
                         in_data[787],
                         in_data[517]
                    }),
            .out_data(lut_275_out)
        );

reg   lut_275_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_275_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_275_ff <= lut_275_out;
    end
end

assign out_data[275] = lut_275_ff;




// LUT : 276

wire lut_276_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111101011111111111010111110111111010011111110),
            .DEVICE(DEVICE)
        )
    i_lut_276
        (
            .in_data({
                         in_data[475],
                         in_data[741],
                         in_data[432],
                         in_data[581],
                         in_data[985],
                         in_data[988]
                    }),
            .out_data(lut_276_out)
        );

reg   lut_276_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_276_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_276_ff <= lut_276_out;
    end
end

assign out_data[276] = lut_276_ff;




// LUT : 277

wire lut_277_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001111101111000000001000011011011111110011111100001111001010),
            .DEVICE(DEVICE)
        )
    i_lut_277
        (
            .in_data({
                         in_data[249],
                         in_data[598],
                         in_data[139],
                         in_data[693],
                         in_data[371],
                         in_data[86]
                    }),
            .out_data(lut_277_out)
        );

reg   lut_277_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_277_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_277_ff <= lut_277_out;
    end
end

assign out_data[277] = lut_277_ff;




// LUT : 278

wire lut_278_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110110101011000000000000001010111111101010110000111000000010),
            .DEVICE(DEVICE)
        )
    i_lut_278
        (
            .in_data({
                         in_data[266],
                         in_data[616],
                         in_data[672],
                         in_data[967],
                         in_data[258],
                         in_data[70]
                    }),
            .out_data(lut_278_out)
        );

reg   lut_278_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_278_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_278_ff <= lut_278_out;
    end
end

assign out_data[278] = lut_278_ff;




// LUT : 279

wire lut_279_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000001010110000100010001010000010101000101010001000101010101000),
            .DEVICE(DEVICE)
        )
    i_lut_279
        (
            .in_data({
                         in_data[941],
                         in_data[650],
                         in_data[135],
                         in_data[845],
                         in_data[306],
                         in_data[448]
                    }),
            .out_data(lut_279_out)
        );

reg   lut_279_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_279_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_279_ff <= lut_279_out;
    end
end

assign out_data[279] = lut_279_ff;




// LUT : 280

wire lut_280_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010100110000010100110100001001110110111111101101010011100110),
            .DEVICE(DEVICE)
        )
    i_lut_280
        (
            .in_data({
                         in_data[806],
                         in_data[396],
                         in_data[600],
                         in_data[7],
                         in_data[452],
                         in_data[781]
                    }),
            .out_data(lut_280_out)
        );

reg   lut_280_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_280_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_280_ff <= lut_280_out;
    end
end

assign out_data[280] = lut_280_ff;




// LUT : 281

wire lut_281_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100000001000000010001010101000000000000000000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_281
        (
            .in_data({
                         in_data[545],
                         in_data[164],
                         in_data[898],
                         in_data[437],
                         in_data[129],
                         in_data[906]
                    }),
            .out_data(lut_281_out)
        );

reg   lut_281_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_281_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_281_ff <= lut_281_out;
    end
end

assign out_data[281] = lut_281_ff;




// LUT : 282

wire lut_282_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110011001000000000000101010011111000111110000001000001010000),
            .DEVICE(DEVICE)
        )
    i_lut_282
        (
            .in_data({
                         in_data[274],
                         in_data[238],
                         in_data[181],
                         in_data[843],
                         in_data[972],
                         in_data[264]
                    }),
            .out_data(lut_282_out)
        );

reg   lut_282_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_282_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_282_ff <= lut_282_out;
    end
end

assign out_data[282] = lut_282_ff;




// LUT : 283

wire lut_283_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111100101111000011000000000011101110110001011110110011000101),
            .DEVICE(DEVICE)
        )
    i_lut_283
        (
            .in_data({
                         in_data[101],
                         in_data[425],
                         in_data[443],
                         in_data[1],
                         in_data[207],
                         in_data[654]
                    }),
            .out_data(lut_283_out)
        );

reg   lut_283_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_283_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_283_ff <= lut_283_out;
    end
end

assign out_data[283] = lut_283_ff;




// LUT : 284

wire lut_284_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111111111111011100111111111110111111111111110011001101111111),
            .DEVICE(DEVICE)
        )
    i_lut_284
        (
            .in_data({
                         in_data[27],
                         in_data[971],
                         in_data[931],
                         in_data[154],
                         in_data[996],
                         in_data[900]
                    }),
            .out_data(lut_284_out)
        );

reg   lut_284_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_284_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_284_ff <= lut_284_out;
    end
end

assign out_data[284] = lut_284_ff;




// LUT : 285

wire lut_285_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111101111110011111100111101001111110011110100111111001111),
            .DEVICE(DEVICE)
        )
    i_lut_285
        (
            .in_data({
                         in_data[667],
                         in_data[549],
                         in_data[669],
                         in_data[877],
                         in_data[839],
                         in_data[605]
                    }),
            .out_data(lut_285_out)
        );

reg   lut_285_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_285_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_285_ff <= lut_285_out;
    end
end

assign out_data[285] = lut_285_ff;




// LUT : 286

wire lut_286_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000001011111010100000101111111101010111111111101000011111111),
            .DEVICE(DEVICE)
        )
    i_lut_286
        (
            .in_data({
                         in_data[764],
                         in_data[547],
                         in_data[151],
                         in_data[758],
                         in_data[237],
                         in_data[921]
                    }),
            .out_data(lut_286_out)
        );

reg   lut_286_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_286_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_286_ff <= lut_286_out;
    end
end

assign out_data[286] = lut_286_ff;




// LUT : 287

wire lut_287_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000011010101111111111111110111110000111011111111110011111111),
            .DEVICE(DEVICE)
        )
    i_lut_287
        (
            .in_data({
                         in_data[610],
                         in_data[1002],
                         in_data[889],
                         in_data[1013],
                         in_data[982],
                         in_data[459]
                    }),
            .out_data(lut_287_out)
        );

reg   lut_287_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_287_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_287_ff <= lut_287_out;
    end
end

assign out_data[287] = lut_287_ff;




// LUT : 288

wire lut_288_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100000000101100010000000000000000001001001001010010010100101),
            .DEVICE(DEVICE)
        )
    i_lut_288
        (
            .in_data({
                         in_data[762],
                         in_data[287],
                         in_data[378],
                         in_data[201],
                         in_data[797],
                         in_data[848]
                    }),
            .out_data(lut_288_out)
        );

reg   lut_288_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_288_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_288_ff <= lut_288_out;
    end
end

assign out_data[288] = lut_288_ff;




// LUT : 289

wire lut_289_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000001000100000000000000000011000101000000010000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_289
        (
            .in_data({
                         in_data[39],
                         in_data[734],
                         in_data[429],
                         in_data[619],
                         in_data[88],
                         in_data[214]
                    }),
            .out_data(lut_289_out)
        );

reg   lut_289_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_289_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_289_ff <= lut_289_out;
    end
end

assign out_data[289] = lut_289_ff;




// LUT : 290

wire lut_290_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111110111111111111100101111101011110000101110001010),
            .DEVICE(DEVICE)
        )
    i_lut_290
        (
            .in_data({
                         in_data[1008],
                         in_data[17],
                         in_data[377],
                         in_data[305],
                         in_data[481],
                         in_data[901]
                    }),
            .out_data(lut_290_out)
        );

reg   lut_290_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_290_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_290_ff <= lut_290_out;
    end
end

assign out_data[290] = lut_290_ff;




// LUT : 291

wire lut_291_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101111111011111111111111111110000110101100001000111111111110000),
            .DEVICE(DEVICE)
        )
    i_lut_291
        (
            .in_data({
                         in_data[634],
                         in_data[844],
                         in_data[413],
                         in_data[957],
                         in_data[89],
                         in_data[1012]
                    }),
            .out_data(lut_291_out)
        );

reg   lut_291_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_291_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_291_ff <= lut_291_out;
    end
end

assign out_data[291] = lut_291_ff;




// LUT : 292

wire lut_292_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011011101011111001110110001001100000000000000000001000100010001),
            .DEVICE(DEVICE)
        )
    i_lut_292
        (
            .in_data({
                         in_data[188],
                         in_data[816],
                         in_data[817],
                         in_data[354],
                         in_data[441],
                         in_data[52]
                    }),
            .out_data(lut_292_out)
        );

reg   lut_292_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_292_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_292_ff <= lut_292_out;
    end
end

assign out_data[292] = lut_292_ff;




// LUT : 293

wire lut_293_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111001111111111111101101000011011110101011111111111111111101),
            .DEVICE(DEVICE)
        )
    i_lut_293
        (
            .in_data({
                         in_data[825],
                         in_data[446],
                         in_data[66],
                         in_data[293],
                         in_data[671],
                         in_data[662]
                    }),
            .out_data(lut_293_out)
        );

reg   lut_293_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_293_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_293_ff <= lut_293_out;
    end
end

assign out_data[293] = lut_293_ff;




// LUT : 294

wire lut_294_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001100000100011000110010010000000011000000111001111110010011100),
            .DEVICE(DEVICE)
        )
    i_lut_294
        (
            .in_data({
                         in_data[586],
                         in_data[861],
                         in_data[866],
                         in_data[158],
                         in_data[576],
                         in_data[965]
                    }),
            .out_data(lut_294_out)
        );

reg   lut_294_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_294_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_294_ff <= lut_294_out;
    end
end

assign out_data[294] = lut_294_ff;




// LUT : 295

wire lut_295_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000100110101111111111111110100010001010101010011110101111111),
            .DEVICE(DEVICE)
        )
    i_lut_295
        (
            .in_data({
                         in_data[614],
                         in_data[822],
                         in_data[709],
                         in_data[310],
                         in_data[580],
                         in_data[449]
                    }),
            .out_data(lut_295_out)
        );

reg   lut_295_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_295_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_295_ff <= lut_295_out;
    end
end

assign out_data[295] = lut_295_ff;




// LUT : 296

wire lut_296_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101111010011101100110000000011111111101100110011101100000000),
            .DEVICE(DEVICE)
        )
    i_lut_296
        (
            .in_data({
                         in_data[955],
                         in_data[885],
                         in_data[570],
                         in_data[681],
                         in_data[728],
                         in_data[608]
                    }),
            .out_data(lut_296_out)
        );

reg   lut_296_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_296_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_296_ff <= lut_296_out;
    end
end

assign out_data[296] = lut_296_ff;




// LUT : 297

wire lut_297_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011101111111011101110111111111110111011111111111011101111111011),
            .DEVICE(DEVICE)
        )
    i_lut_297
        (
            .in_data({
                         in_data[962],
                         in_data[854],
                         in_data[324],
                         in_data[720],
                         in_data[160],
                         in_data[138]
                    }),
            .out_data(lut_297_out)
        );

reg   lut_297_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_297_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_297_ff <= lut_297_out;
    end
end

assign out_data[297] = lut_297_ff;




// LUT : 298

wire lut_298_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110001100111011111111110010111111001111001110101111110000),
            .DEVICE(DEVICE)
        )
    i_lut_298
        (
            .in_data({
                         in_data[45],
                         in_data[578],
                         in_data[93],
                         in_data[84],
                         in_data[56],
                         in_data[259]
                    }),
            .out_data(lut_298_out)
        );

reg   lut_298_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_298_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_298_ff <= lut_298_out;
    end
end

assign out_data[298] = lut_298_ff;




// LUT : 299

wire lut_299_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111011111111010011001111111111101111111111111010110011111100),
            .DEVICE(DEVICE)
        )
    i_lut_299
        (
            .in_data({
                         in_data[442],
                         in_data[11],
                         in_data[384],
                         in_data[611],
                         in_data[785],
                         in_data[940]
                    }),
            .out_data(lut_299_out)
        );

reg   lut_299_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_299_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_299_ff <= lut_299_out;
    end
end

assign out_data[299] = lut_299_ff;




// LUT : 300

wire lut_300_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000001000000100000000100000000000000000000010000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_300
        (
            .in_data({
                         in_data[40],
                         in_data[656],
                         in_data[869],
                         in_data[124],
                         in_data[978],
                         in_data[191]
                    }),
            .out_data(lut_300_out)
        );

reg   lut_300_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_300_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_300_ff <= lut_300_out;
    end
end

assign out_data[300] = lut_300_ff;




// LUT : 301

wire lut_301_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111001111110000100001111011110100010001011100011010101101101),
            .DEVICE(DEVICE)
        )
    i_lut_301
        (
            .in_data({
                         in_data[715],
                         in_data[841],
                         in_data[585],
                         in_data[942],
                         in_data[540],
                         in_data[697]
                    }),
            .out_data(lut_301_out)
        );

reg   lut_301_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_301_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_301_ff <= lut_301_out;
    end
end

assign out_data[301] = lut_301_ff;




// LUT : 302

wire lut_302_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110011001100110011010100110011111111110011111100111111001101),
            .DEVICE(DEVICE)
        )
    i_lut_302
        (
            .in_data({
                         in_data[179],
                         in_data[339],
                         in_data[928],
                         in_data[873],
                         in_data[960],
                         in_data[383]
                    }),
            .out_data(lut_302_out)
        );

reg   lut_302_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_302_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_302_ff <= lut_302_out;
    end
end

assign out_data[302] = lut_302_ff;




// LUT : 303

wire lut_303_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010101010101110000000001100110000111010111111101111111111001111),
            .DEVICE(DEVICE)
        )
    i_lut_303
        (
            .in_data({
                         in_data[914],
                         in_data[327],
                         in_data[224],
                         in_data[766],
                         in_data[61],
                         in_data[595]
                    }),
            .out_data(lut_303_out)
        );

reg   lut_303_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_303_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_303_ff <= lut_303_out;
    end
end

assign out_data[303] = lut_303_ff;




// LUT : 304

wire lut_304_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111111111111000111111111111100001111111111110000111111111101),
            .DEVICE(DEVICE)
        )
    i_lut_304
        (
            .in_data({
                         in_data[879],
                         in_data[945],
                         in_data[769],
                         in_data[23],
                         in_data[171],
                         in_data[999]
                    }),
            .out_data(lut_304_out)
        );

reg   lut_304_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_304_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_304_ff <= lut_304_out;
    end
end

assign out_data[304] = lut_304_ff;




// LUT : 305

wire lut_305_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001111101001101000000000000000000001111000000000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_305
        (
            .in_data({
                         in_data[870],
                         in_data[16],
                         in_data[281],
                         in_data[42],
                         in_data[85],
                         in_data[337]
                    }),
            .out_data(lut_305_out)
        );

reg   lut_305_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_305_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_305_ff <= lut_305_out;
    end
end

assign out_data[305] = lut_305_ff;




// LUT : 306

wire lut_306_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111100101010111111111011101111001110100010001111111100111010),
            .DEVICE(DEVICE)
        )
    i_lut_306
        (
            .in_data({
                         in_data[260],
                         in_data[648],
                         in_data[863],
                         in_data[95],
                         in_data[563],
                         in_data[130]
                    }),
            .out_data(lut_306_out)
        );

reg   lut_306_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_306_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_306_ff <= lut_306_out;
    end
end

assign out_data[306] = lut_306_ff;




// LUT : 307

wire lut_307_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110111110011111001111010111000011001111000100000000010101011),
            .DEVICE(DEVICE)
        )
    i_lut_307
        (
            .in_data({
                         in_data[137],
                         in_data[268],
                         in_data[918],
                         in_data[329],
                         in_data[882],
                         in_data[119]
                    }),
            .out_data(lut_307_out)
        );

reg   lut_307_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_307_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_307_ff <= lut_307_out;
    end
end

assign out_data[307] = lut_307_ff;




// LUT : 308

wire lut_308_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111110101110111111111010111011100000101000001010010010100000),
            .DEVICE(DEVICE)
        )
    i_lut_308
        (
            .in_data({
                         in_data[526],
                         in_data[646],
                         in_data[635],
                         in_data[462],
                         in_data[794],
                         in_data[338]
                    }),
            .out_data(lut_308_out)
        );

reg   lut_308_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_308_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_308_ff <= lut_308_out;
    end
end

assign out_data[308] = lut_308_ff;




// LUT : 309

wire lut_309_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001000000000001000100000000000100010000000100010101100001010),
            .DEVICE(DEVICE)
        )
    i_lut_309
        (
            .in_data({
                         in_data[363],
                         in_data[779],
                         in_data[742],
                         in_data[195],
                         in_data[814],
                         in_data[350]
                    }),
            .out_data(lut_309_out)
        );

reg   lut_309_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_309_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_309_ff <= lut_309_out;
    end
end

assign out_data[309] = lut_309_ff;




// LUT : 310

wire lut_310_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000011110100000000000100000000100011001000001111001111111111),
            .DEVICE(DEVICE)
        )
    i_lut_310
        (
            .in_data({
                         in_data[707],
                         in_data[621],
                         in_data[239],
                         in_data[891],
                         in_data[473],
                         in_data[18]
                    }),
            .out_data(lut_310_out)
        );

reg   lut_310_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_310_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_310_ff <= lut_310_out;
    end
end

assign out_data[310] = lut_310_ff;




// LUT : 311

wire lut_311_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100010011110100010000000100000001000100111101011100010011000000),
            .DEVICE(DEVICE)
        )
    i_lut_311
        (
            .in_data({
                         in_data[405],
                         in_data[122],
                         in_data[796],
                         in_data[166],
                         in_data[63],
                         in_data[412]
                    }),
            .out_data(lut_311_out)
        );

reg   lut_311_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_311_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_311_ff <= lut_311_out;
    end
end

assign out_data[311] = lut_311_ff;




// LUT : 312

wire lut_312_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111011111111111111111111111111111010101011111111),
            .DEVICE(DEVICE)
        )
    i_lut_312
        (
            .in_data({
                         in_data[793],
                         in_data[87],
                         in_data[620],
                         in_data[874],
                         in_data[468],
                         in_data[491]
                    }),
            .out_data(lut_312_out)
        );

reg   lut_312_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_312_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_312_ff <= lut_312_out;
    end
end

assign out_data[312] = lut_312_ff;




// LUT : 313

wire lut_313_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100110000001110110111011000110111011100100111001101100000011),
            .DEVICE(DEVICE)
        )
    i_lut_313
        (
            .in_data({
                         in_data[91],
                         in_data[34],
                         in_data[444],
                         in_data[271],
                         in_data[190],
                         in_data[262]
                    }),
            .out_data(lut_313_out)
        );

reg   lut_313_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_313_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_313_ff <= lut_313_out;
    end
end

assign out_data[313] = lut_313_ff;




// LUT : 314

wire lut_314_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111011111110011111111101010111110110111111000111111),
            .DEVICE(DEVICE)
        )
    i_lut_314
        (
            .in_data({
                         in_data[744],
                         in_data[120],
                         in_data[353],
                         in_data[831],
                         in_data[289],
                         in_data[790]
                    }),
            .out_data(lut_314_out)
        );

reg   lut_314_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_314_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_314_ff <= lut_314_out;
    end
end

assign out_data[314] = lut_314_ff;




// LUT : 315

wire lut_315_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010000000100110000001011010001000010001111110110101010111111111),
            .DEVICE(DEVICE)
        )
    i_lut_315
        (
            .in_data({
                         in_data[977],
                         in_data[474],
                         in_data[435],
                         in_data[389],
                         in_data[640],
                         in_data[772]
                    }),
            .out_data(lut_315_out)
        );

reg   lut_315_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_315_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_315_ff <= lut_315_out;
    end
end

assign out_data[315] = lut_315_ff;




// LUT : 316

wire lut_316_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010000000100000000000001010000000001101000001110000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_316
        (
            .in_data({
                         in_data[857],
                         in_data[632],
                         in_data[926],
                         in_data[663],
                         in_data[317],
                         in_data[1023]
                    }),
            .out_data(lut_316_out)
        );

reg   lut_316_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_316_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_316_ff <= lut_316_out;
    end
end

assign out_data[316] = lut_316_ff;




// LUT : 317

wire lut_317_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0110111111111111111111101111111110001111001111111100100010101011),
            .DEVICE(DEVICE)
        )
    i_lut_317
        (
            .in_data({
                         in_data[2],
                         in_data[351],
                         in_data[688],
                         in_data[54],
                         in_data[250],
                         in_data[603]
                    }),
            .out_data(lut_317_out)
        );

reg   lut_317_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_317_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_317_ff <= lut_317_out;
    end
end

assign out_data[317] = lut_317_ff;




// LUT : 318

wire lut_318_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010011111111111100001111111111110000111111111101000011111111),
            .DEVICE(DEVICE)
        )
    i_lut_318
        (
            .in_data({
                         in_data[267],
                         in_data[735],
                         in_data[193],
                         in_data[551],
                         in_data[460],
                         in_data[370]
                    }),
            .out_data(lut_318_out)
        );

reg   lut_318_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_318_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_318_ff <= lut_318_out;
    end
end

assign out_data[318] = lut_318_ff;




// LUT : 319

wire lut_319_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000001010111011101000101001001100000010001110100010001100),
            .DEVICE(DEVICE)
        )
    i_lut_319
        (
            .in_data({
                         in_data[323],
                         in_data[424],
                         in_data[647],
                         in_data[930],
                         in_data[465],
                         in_data[205]
                    }),
            .out_data(lut_319_out)
        );

reg   lut_319_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_319_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_319_ff <= lut_319_out;
    end
end

assign out_data[319] = lut_319_ff;




// LUT : 320

wire lut_320_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001001000000000000100110000110011001000100000000000000100),
            .DEVICE(DEVICE)
        )
    i_lut_320
        (
            .in_data({
                         in_data[187],
                         in_data[864],
                         in_data[172],
                         in_data[229],
                         in_data[823],
                         in_data[208]
                    }),
            .out_data(lut_320_out)
        );

reg   lut_320_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_320_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_320_ff <= lut_320_out;
    end
end

assign out_data[320] = lut_320_ff;




// LUT : 321

wire lut_321_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111000000000101011101100001110101110111011101111111011001101),
            .DEVICE(DEVICE)
        )
    i_lut_321
        (
            .in_data({
                         in_data[986],
                         in_data[6],
                         in_data[265],
                         in_data[835],
                         in_data[157],
                         in_data[77]
                    }),
            .out_data(lut_321_out)
        );

reg   lut_321_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_321_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_321_ff <= lut_321_out;
    end
end

assign out_data[321] = lut_321_ff;




// LUT : 322

wire lut_322_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000000111001100110101110000111111111111110001001111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_322
        (
            .in_data({
                         in_data[313],
                         in_data[664],
                         in_data[630],
                         in_data[415],
                         in_data[498],
                         in_data[602]
                    }),
            .out_data(lut_322_out)
        );

reg   lut_322_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_322_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_322_ff <= lut_322_out;
    end
end

assign out_data[322] = lut_322_ff;




// LUT : 323

wire lut_323_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000001111000000000000000011001110000011111100110000101011),
            .DEVICE(DEVICE)
        )
    i_lut_323
        (
            .in_data({
                         in_data[357],
                         in_data[434],
                         in_data[231],
                         in_data[704],
                         in_data[393],
                         in_data[567]
                    }),
            .out_data(lut_323_out)
        );

reg   lut_323_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_323_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_323_ff <= lut_323_out;
    end
end

assign out_data[323] = lut_323_ff;




// LUT : 324

wire lut_324_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111110100111101100000010111101001011100000111101101101101011),
            .DEVICE(DEVICE)
        )
    i_lut_324
        (
            .in_data({
                         in_data[725],
                         in_data[893],
                         in_data[763],
                         in_data[326],
                         in_data[24],
                         in_data[653]
                    }),
            .out_data(lut_324_out)
        );

reg   lut_324_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_324_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_324_ff <= lut_324_out;
    end
end

assign out_data[324] = lut_324_ff;




// LUT : 325

wire lut_325_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000001110000000000000000000000000000111100000000),
            .DEVICE(DEVICE)
        )
    i_lut_325
        (
            .in_data({
                         in_data[1003],
                         in_data[394],
                         in_data[1011],
                         in_data[445],
                         in_data[270],
                         in_data[850]
                    }),
            .out_data(lut_325_out)
        );

reg   lut_325_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_325_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_325_ff <= lut_325_out;
    end
end

assign out_data[325] = lut_325_ff;




// LUT : 326

wire lut_326_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001100100001000000010000000000000000000000000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_326
        (
            .in_data({
                         in_data[561],
                         in_data[564],
                         in_data[624],
                         in_data[542],
                         in_data[519],
                         in_data[736]
                    }),
            .out_data(lut_326_out)
        );

reg   lut_326_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_326_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_326_ff <= lut_326_out;
    end
end

assign out_data[326] = lut_326_ff;




// LUT : 327

wire lut_327_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000010011000000000000000000000101001000100101010111001000),
            .DEVICE(DEVICE)
        )
    i_lut_327
        (
            .in_data({
                         in_data[811],
                         in_data[272],
                         in_data[686],
                         in_data[538],
                         in_data[499],
                         in_data[103]
                    }),
            .out_data(lut_327_out)
        );

reg   lut_327_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_327_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_327_ff <= lut_327_out;
    end
end

assign out_data[327] = lut_327_ff;




// LUT : 328

wire lut_328_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011001111111111111111101001101011111111111111101111111111111010),
            .DEVICE(DEVICE)
        )
    i_lut_328
        (
            .in_data({
                         in_data[116],
                         in_data[810],
                         in_data[275],
                         in_data[248],
                         in_data[430],
                         in_data[153]
                    }),
            .out_data(lut_328_out)
        );

reg   lut_328_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_328_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_328_ff <= lut_328_out;
    end
end

assign out_data[328] = lut_328_ff;




// LUT : 329

wire lut_329_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101011001010011111111011111110011101001010001001111101001100101),
            .DEVICE(DEVICE)
        )
    i_lut_329
        (
            .in_data({
                         in_data[699],
                         in_data[859],
                         in_data[60],
                         in_data[767],
                         in_data[471],
                         in_data[680]
                    }),
            .out_data(lut_329_out)
        );

reg   lut_329_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_329_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_329_ff <= lut_329_out;
    end
end

assign out_data[329] = lut_329_ff;




// LUT : 330

wire lut_330_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111111111111000101010001000111111111100011001111001100000001),
            .DEVICE(DEVICE)
        )
    i_lut_330
        (
            .in_data({
                         in_data[760],
                         in_data[949],
                         in_data[69],
                         in_data[902],
                         in_data[32],
                         in_data[283]
                    }),
            .out_data(lut_330_out)
        );

reg   lut_330_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_330_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_330_ff <= lut_330_out;
    end
end

assign out_data[330] = lut_330_ff;




// LUT : 331

wire lut_331_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100010010001001100101001111110001000000100010000000000010001000),
            .DEVICE(DEVICE)
        )
    i_lut_331
        (
            .in_data({
                         in_data[636],
                         in_data[209],
                         in_data[748],
                         in_data[131],
                         in_data[912],
                         in_data[661]
                    }),
            .out_data(lut_331_out)
        );

reg   lut_331_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_331_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_331_ff <= lut_331_out;
    end
end

assign out_data[331] = lut_331_ff;




// LUT : 332

wire lut_332_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101111111011011001101111110110111011101110111010111101011011),
            .DEVICE(DEVICE)
        )
    i_lut_332
        (
            .in_data({
                         in_data[504],
                         in_data[537],
                         in_data[246],
                         in_data[476],
                         in_data[995],
                         in_data[502]
                    }),
            .out_data(lut_332_out)
        );

reg   lut_332_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_332_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_332_ff <= lut_332_out;
    end
end

assign out_data[332] = lut_332_ff;




// LUT : 333

wire lut_333_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000000000000000110010000011111000000000001010),
            .DEVICE(DEVICE)
        )
    i_lut_333
        (
            .in_data({
                         in_data[513],
                         in_data[539],
                         in_data[484],
                         in_data[652],
                         in_data[269],
                         in_data[182]
                    }),
            .out_data(lut_333_out)
        );

reg   lut_333_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_333_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_333_ff <= lut_333_out;
    end
end

assign out_data[333] = lut_333_ff;




// LUT : 334

wire lut_334_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101100010011111111111011111111111111111111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_334
        (
            .in_data({
                         in_data[573],
                         in_data[406],
                         in_data[802],
                         in_data[968],
                         in_data[792],
                         in_data[387]
                    }),
            .out_data(lut_334_out)
        );

reg   lut_334_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_334_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_334_ff <= lut_334_out;
    end
end

assign out_data[334] = lut_334_ff;




// LUT : 335

wire lut_335_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100010110000110010001111111111111010101100001111001011110100),
            .DEVICE(DEVICE)
        )
    i_lut_335
        (
            .in_data({
                         in_data[756],
                         in_data[302],
                         in_data[490],
                         in_data[950],
                         in_data[447],
                         in_data[251]
                    }),
            .out_data(lut_335_out)
        );

reg   lut_335_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_335_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_335_ff <= lut_335_out;
    end
end

assign out_data[335] = lut_335_ff;




// LUT : 336

wire lut_336_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000101001011101101111110111100011111111111010101111111111010001),
            .DEVICE(DEVICE)
        )
    i_lut_336
        (
            .in_data({
                         in_data[64],
                         in_data[399],
                         in_data[903],
                         in_data[932],
                         in_data[613],
                         in_data[73]
                    }),
            .out_data(lut_336_out)
        );

reg   lut_336_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_336_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_336_ff <= lut_336_out;
    end
end

assign out_data[336] = lut_336_ff;




// LUT : 337

wire lut_337_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110001110000010001010001000101011101000100000000010100000001),
            .DEVICE(DEVICE)
        )
    i_lut_337
        (
            .in_data({
                         in_data[981],
                         in_data[192],
                         in_data[28],
                         in_data[544],
                         in_data[176],
                         in_data[703]
                    }),
            .out_data(lut_337_out)
        );

reg   lut_337_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_337_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_337_ff <= lut_337_out;
    end
end

assign out_data[337] = lut_337_ff;




// LUT : 338

wire lut_338_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000011110000011100010101000100000000000001010100010100001100),
            .DEVICE(DEVICE)
        )
    i_lut_338
        (
            .in_data({
                         in_data[366],
                         in_data[334],
                         in_data[202],
                         in_data[152],
                         in_data[303],
                         in_data[106]
                    }),
            .out_data(lut_338_out)
        );

reg   lut_338_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_338_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_338_ff <= lut_338_out;
    end
end

assign out_data[338] = lut_338_ff;




// LUT : 339

wire lut_339_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010000000100111101000000011100000000000000001100010100000101),
            .DEVICE(DEVICE)
        )
    i_lut_339
        (
            .in_data({
                         in_data[165],
                         in_data[974],
                         in_data[245],
                         in_data[358],
                         in_data[917],
                         in_data[9]
                    }),
            .out_data(lut_339_out)
        );

reg   lut_339_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_339_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_339_ff <= lut_339_out;
    end
end

assign out_data[339] = lut_339_ff;




// LUT : 340

wire lut_340_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111101011111111111101101101011011111110111111100110001011111),
            .DEVICE(DEVICE)
        )
    i_lut_340
        (
            .in_data({
                         in_data[974],
                         in_data[385],
                         in_data[360],
                         in_data[288],
                         in_data[486],
                         in_data[702]
                    }),
            .out_data(lut_340_out)
        );

reg   lut_340_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_340_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_340_ff <= lut_340_out;
    end
end

assign out_data[340] = lut_340_ff;




// LUT : 341

wire lut_341_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100000011001000110011001100011000000110000011110000000011000101),
            .DEVICE(DEVICE)
        )
    i_lut_341
        (
            .in_data({
                         in_data[64],
                         in_data[55],
                         in_data[10],
                         in_data[275],
                         in_data[161],
                         in_data[303]
                    }),
            .out_data(lut_341_out)
        );

reg   lut_341_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_341_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_341_ff <= lut_341_out;
    end
end

assign out_data[341] = lut_341_ff;




// LUT : 342

wire lut_342_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010001100010000111111110000100111111111000100001110111101001100),
            .DEVICE(DEVICE)
        )
    i_lut_342
        (
            .in_data({
                         in_data[59],
                         in_data[345],
                         in_data[895],
                         in_data[580],
                         in_data[711],
                         in_data[322]
                    }),
            .out_data(lut_342_out)
        );

reg   lut_342_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_342_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_342_ff <= lut_342_out;
    end
end

assign out_data[342] = lut_342_ff;




// LUT : 343

wire lut_343_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110001111110010001011111111111100000010111100100000111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_343
        (
            .in_data({
                         in_data[599],
                         in_data[289],
                         in_data[866],
                         in_data[617],
                         in_data[590],
                         in_data[713]
                    }),
            .out_data(lut_343_out)
        );

reg   lut_343_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_343_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_343_ff <= lut_343_out;
    end
end

assign out_data[343] = lut_343_ff;




// LUT : 344

wire lut_344_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110011101100111001001111110000000000110000000000000011000000),
            .DEVICE(DEVICE)
        )
    i_lut_344
        (
            .in_data({
                         in_data[5],
                         in_data[210],
                         in_data[127],
                         in_data[319],
                         in_data[133],
                         in_data[148]
                    }),
            .out_data(lut_344_out)
        );

reg   lut_344_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_344_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_344_ff <= lut_344_out;
    end
end

assign out_data[344] = lut_344_ff;




// LUT : 345

wire lut_345_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111101110111111111110101111101110111000000000100011100000000),
            .DEVICE(DEVICE)
        )
    i_lut_345
        (
            .in_data({
                         in_data[65],
                         in_data[605],
                         in_data[164],
                         in_data[1022],
                         in_data[9],
                         in_data[744]
                    }),
            .out_data(lut_345_out)
        );

reg   lut_345_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_345_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_345_ff <= lut_345_out;
    end
end

assign out_data[345] = lut_345_ff;




// LUT : 346

wire lut_346_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000101010101001101111111111111111111111111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_346
        (
            .in_data({
                         in_data[477],
                         in_data[571],
                         in_data[48],
                         in_data[588],
                         in_data[682],
                         in_data[812]
                    }),
            .out_data(lut_346_out)
        );

reg   lut_346_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_346_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_346_ff <= lut_346_out;
    end
end

assign out_data[346] = lut_346_ff;




// LUT : 347

wire lut_347_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000001010000000001000101000001100000010001100111000001010),
            .DEVICE(DEVICE)
        )
    i_lut_347
        (
            .in_data({
                         in_data[634],
                         in_data[969],
                         in_data[863],
                         in_data[338],
                         in_data[459],
                         in_data[261]
                    }),
            .out_data(lut_347_out)
        );

reg   lut_347_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_347_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_347_ff <= lut_347_out;
    end
end

assign out_data[347] = lut_347_ff;




// LUT : 348

wire lut_348_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001100101010111111111010110000101011001101111010111111101110),
            .DEVICE(DEVICE)
        )
    i_lut_348
        (
            .in_data({
                         in_data[19],
                         in_data[805],
                         in_data[245],
                         in_data[779],
                         in_data[260],
                         in_data[92]
                    }),
            .out_data(lut_348_out)
        );

reg   lut_348_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_348_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_348_ff <= lut_348_out;
    end
end

assign out_data[348] = lut_348_ff;




// LUT : 349

wire lut_349_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000000110000000000000000000011010000110101000100000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_349
        (
            .in_data({
                         in_data[388],
                         in_data[623],
                         in_data[649],
                         in_data[918],
                         in_data[359],
                         in_data[873]
                    }),
            .out_data(lut_349_out)
        );

reg   lut_349_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_349_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_349_ff <= lut_349_out;
    end
end

assign out_data[349] = lut_349_ff;




// LUT : 350

wire lut_350_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101000000011011110110101000000001000000000100111000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_350
        (
            .in_data({
                         in_data[379],
                         in_data[87],
                         in_data[225],
                         in_data[71],
                         in_data[405],
                         in_data[633]
                    }),
            .out_data(lut_350_out)
        );

reg   lut_350_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_350_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_350_ff <= lut_350_out;
    end
end

assign out_data[350] = lut_350_ff;




// LUT : 351

wire lut_351_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111110111111000000111010111111111111000110100100111100101010),
            .DEVICE(DEVICE)
        )
    i_lut_351
        (
            .in_data({
                         in_data[306],
                         in_data[788],
                         in_data[500],
                         in_data[103],
                         in_data[499],
                         in_data[476]
                    }),
            .out_data(lut_351_out)
        );

reg   lut_351_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_351_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_351_ff <= lut_351_out;
    end
end

assign out_data[351] = lut_351_ff;




// LUT : 352

wire lut_352_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100100000100101100010000000001000000000011001010000000000110000),
            .DEVICE(DEVICE)
        )
    i_lut_352
        (
            .in_data({
                         in_data[657],
                         in_data[496],
                         in_data[201],
                         in_data[931],
                         in_data[731],
                         in_data[554]
                    }),
            .out_data(lut_352_out)
        );

reg   lut_352_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_352_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_352_ff <= lut_352_out;
    end
end

assign out_data[352] = lut_352_ff;




// LUT : 353

wire lut_353_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011101100101011111110111111111111101101111111111100111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_353
        (
            .in_data({
                         in_data[818],
                         in_data[540],
                         in_data[29],
                         in_data[615],
                         in_data[772],
                         in_data[240]
                    }),
            .out_data(lut_353_out)
        );

reg   lut_353_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_353_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_353_ff <= lut_353_out;
    end
end

assign out_data[353] = lut_353_ff;




// LUT : 354

wire lut_354_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111110111011111110111111111111111111101111101010000),
            .DEVICE(DEVICE)
        )
    i_lut_354
        (
            .in_data({
                         in_data[773],
                         in_data[608],
                         in_data[390],
                         in_data[628],
                         in_data[665],
                         in_data[233]
                    }),
            .out_data(lut_354_out)
        );

reg   lut_354_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_354_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_354_ff <= lut_354_out;
    end
end

assign out_data[354] = lut_354_ff;




// LUT : 355

wire lut_355_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000001111111111101110101011110000010011101101111010101010111111),
            .DEVICE(DEVICE)
        )
    i_lut_355
        (
            .in_data({
                         in_data[977],
                         in_data[544],
                         in_data[998],
                         in_data[159],
                         in_data[515],
                         in_data[817]
                    }),
            .out_data(lut_355_out)
        );

reg   lut_355_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_355_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_355_ff <= lut_355_out;
    end
end

assign out_data[355] = lut_355_ff;




// LUT : 356

wire lut_356_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001111110000111001111100010000100111111011011000111111101100),
            .DEVICE(DEVICE)
        )
    i_lut_356
        (
            .in_data({
                         in_data[171],
                         in_data[453],
                         in_data[901],
                         in_data[28],
                         in_data[869],
                         in_data[920]
                    }),
            .out_data(lut_356_out)
        );

reg   lut_356_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_356_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_356_ff <= lut_356_out;
    end
end

assign out_data[356] = lut_356_ff;




// LUT : 357

wire lut_357_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110111101101111001001110010111111111111111111110111111101111),
            .DEVICE(DEVICE)
        )
    i_lut_357
        (
            .in_data({
                         in_data[157],
                         in_data[567],
                         in_data[842],
                         in_data[450],
                         in_data[172],
                         in_data[865]
                    }),
            .out_data(lut_357_out)
        );

reg   lut_357_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_357_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_357_ff <= lut_357_out;
    end
end

assign out_data[357] = lut_357_ff;




// LUT : 358

wire lut_358_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101000100000000001101010000000011111111000000000101010100000000),
            .DEVICE(DEVICE)
        )
    i_lut_358
        (
            .in_data({
                         in_data[274],
                         in_data[517],
                         in_data[158],
                         in_data[286],
                         in_data[785],
                         in_data[119]
                    }),
            .out_data(lut_358_out)
        );

reg   lut_358_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_358_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_358_ff <= lut_358_out;
    end
end

assign out_data[358] = lut_358_ff;




// LUT : 359

wire lut_359_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111100001000001011111010101010101010000000000000010000000000),
            .DEVICE(DEVICE)
        )
    i_lut_359
        (
            .in_data({
                         in_data[340],
                         in_data[346],
                         in_data[409],
                         in_data[263],
                         in_data[935],
                         in_data[72]
                    }),
            .out_data(lut_359_out)
        );

reg   lut_359_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_359_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_359_ff <= lut_359_out;
    end
end

assign out_data[359] = lut_359_ff;



endmodule



module MnistStochasticLut6Mlp_sub2
        #(
            parameter DEVICE = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [359:0]  in_data,
            output wire [59:0]  out_data
        );


// LUT : 0

wire lut_0_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010101010000011100010111000001010101000000000111000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_0
        (
            .in_data({
                         in_data[111],
                         in_data[82],
                         in_data[280],
                         in_data[316],
                         in_data[302],
                         in_data[8]
                    }),
            .out_data(lut_0_out)
        );

reg   lut_0_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_0_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_0_ff <= lut_0_out;
    end
end

assign out_data[0] = lut_0_ff;




// LUT : 1

wire lut_1_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111000100110000000100000011000001110111111100110011000101110111),
            .DEVICE(DEVICE)
        )
    i_lut_1
        (
            .in_data({
                         in_data[20],
                         in_data[289],
                         in_data[203],
                         in_data[344],
                         in_data[191],
                         in_data[73]
                    }),
            .out_data(lut_1_out)
        );

reg   lut_1_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1_ff <= lut_1_out;
    end
end

assign out_data[1] = lut_1_ff;




// LUT : 2

wire lut_2_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000011110001000000000111000101110011111111110011000011110111),
            .DEVICE(DEVICE)
        )
    i_lut_2
        (
            .in_data({
                         in_data[310],
                         in_data[148],
                         in_data[47],
                         in_data[10],
                         in_data[278],
                         in_data[71]
                    }),
            .out_data(lut_2_out)
        );

reg   lut_2_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_2_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_2_ff <= lut_2_out;
    end
end

assign out_data[2] = lut_2_ff;




// LUT : 3

wire lut_3_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100000000000101011110000010010001110000010001111111111101111),
            .DEVICE(DEVICE)
        )
    i_lut_3
        (
            .in_data({
                         in_data[330],
                         in_data[120],
                         in_data[98],
                         in_data[178],
                         in_data[44],
                         in_data[133]
                    }),
            .out_data(lut_3_out)
        );

reg   lut_3_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_3_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_3_ff <= lut_3_out;
    end
end

assign out_data[3] = lut_3_ff;




// LUT : 4

wire lut_4_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101111111111001000000011001111111011111111111010000000110011),
            .DEVICE(DEVICE)
        )
    i_lut_4
        (
            .in_data({
                         in_data[132],
                         in_data[234],
                         in_data[48],
                         in_data[129],
                         in_data[259],
                         in_data[334]
                    }),
            .out_data(lut_4_out)
        );

reg   lut_4_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_4_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_4_ff <= lut_4_out;
    end
end

assign out_data[4] = lut_4_ff;




// LUT : 5

wire lut_5_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000000000000000010111000100010000100100000000),
            .DEVICE(DEVICE)
        )
    i_lut_5
        (
            .in_data({
                         in_data[0],
                         in_data[65],
                         in_data[30],
                         in_data[193],
                         in_data[298],
                         in_data[41]
                    }),
            .out_data(lut_5_out)
        );

reg   lut_5_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_5_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_5_ff <= lut_5_out;
    end
end

assign out_data[5] = lut_5_ff;




// LUT : 6

wire lut_6_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000100000001000000010000000000010011000000110001001100000001),
            .DEVICE(DEVICE)
        )
    i_lut_6
        (
            .in_data({
                         in_data[206],
                         in_data[359],
                         in_data[347],
                         in_data[40],
                         in_data[135],
                         in_data[205]
                    }),
            .out_data(lut_6_out)
        );

reg   lut_6_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_6_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_6_ff <= lut_6_out;
    end
end

assign out_data[6] = lut_6_ff;




// LUT : 7

wire lut_7_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010000011111000111110011111101111111111111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_7
        (
            .in_data({
                         in_data[338],
                         in_data[341],
                         in_data[61],
                         in_data[254],
                         in_data[320],
                         in_data[275]
                    }),
            .out_data(lut_7_out)
        );

reg   lut_7_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_7_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_7_ff <= lut_7_out;
    end
end

assign out_data[7] = lut_7_ff;




// LUT : 8

wire lut_8_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101111111111111010111010101010111111111111111111101111101011111),
            .DEVICE(DEVICE)
        )
    i_lut_8
        (
            .in_data({
                         in_data[200],
                         in_data[101],
                         in_data[194],
                         in_data[274],
                         in_data[78],
                         in_data[329]
                    }),
            .out_data(lut_8_out)
        );

reg   lut_8_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_8_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_8_ff <= lut_8_out;
    end
end

assign out_data[8] = lut_8_ff;




// LUT : 9

wire lut_9_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000001101000000000000010000001100000011110100),
            .DEVICE(DEVICE)
        )
    i_lut_9
        (
            .in_data({
                         in_data[157],
                         in_data[322],
                         in_data[265],
                         in_data[327],
                         in_data[141],
                         in_data[355]
                    }),
            .out_data(lut_9_out)
        );

reg   lut_9_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_9_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_9_ff <= lut_9_out;
    end
end

assign out_data[9] = lut_9_ff;




// LUT : 10

wire lut_10_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111110101010100010011010000010001010000010000000100000000000100),
            .DEVICE(DEVICE)
        )
    i_lut_10
        (
            .in_data({
                         in_data[218],
                         in_data[235],
                         in_data[252],
                         in_data[37],
                         in_data[36],
                         in_data[296]
                    }),
            .out_data(lut_10_out)
        );

reg   lut_10_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_10_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_10_ff <= lut_10_out;
    end
end

assign out_data[10] = lut_10_ff;




// LUT : 11

wire lut_11_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101000000000000000000000000000011011101010000001100010000000000),
            .DEVICE(DEVICE)
        )
    i_lut_11
        (
            .in_data({
                         in_data[125],
                         in_data[159],
                         in_data[124],
                         in_data[32],
                         in_data[53],
                         in_data[224]
                    }),
            .out_data(lut_11_out)
        );

reg   lut_11_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_11_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_11_ff <= lut_11_out;
    end
end

assign out_data[11] = lut_11_ff;




// LUT : 12

wire lut_12_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111101111111000101110001000111111111111111110111111100010001),
            .DEVICE(DEVICE)
        )
    i_lut_12
        (
            .in_data({
                         in_data[123],
                         in_data[147],
                         in_data[340],
                         in_data[115],
                         in_data[171],
                         in_data[96]
                    }),
            .out_data(lut_12_out)
        );

reg   lut_12_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_12_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_12_ff <= lut_12_out;
    end
end

assign out_data[12] = lut_12_ff;




// LUT : 13

wire lut_13_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011111111111111000011110011111111111111111100111110111001100011),
            .DEVICE(DEVICE)
        )
    i_lut_13
        (
            .in_data({
                         in_data[181],
                         in_data[222],
                         in_data[263],
                         in_data[168],
                         in_data[128],
                         in_data[232]
                    }),
            .out_data(lut_13_out)
        );

reg   lut_13_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_13_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_13_ff <= lut_13_out;
    end
end

assign out_data[13] = lut_13_ff;




// LUT : 14

wire lut_14_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000100000000000000000000000000010111100000010),
            .DEVICE(DEVICE)
        )
    i_lut_14
        (
            .in_data({
                         in_data[293],
                         in_data[276],
                         in_data[352],
                         in_data[104],
                         in_data[19],
                         in_data[94]
                    }),
            .out_data(lut_14_out)
        );

reg   lut_14_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_14_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_14_ff <= lut_14_out;
    end
end

assign out_data[14] = lut_14_ff;




// LUT : 15

wire lut_15_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100111111111111110111111111111111001101111111111101111111011111),
            .DEVICE(DEVICE)
        )
    i_lut_15
        (
            .in_data({
                         in_data[144],
                         in_data[79],
                         in_data[267],
                         in_data[272],
                         in_data[317],
                         in_data[112]
                    }),
            .out_data(lut_15_out)
        );

reg   lut_15_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_15_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_15_ff <= lut_15_out;
    end
end

assign out_data[15] = lut_15_ff;




// LUT : 16

wire lut_16_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111011111111111011111111111100001000110011000010111011101111),
            .DEVICE(DEVICE)
        )
    i_lut_16
        (
            .in_data({
                         in_data[353],
                         in_data[116],
                         in_data[337],
                         in_data[58],
                         in_data[97],
                         in_data[247]
                    }),
            .out_data(lut_16_out)
        );

reg   lut_16_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_16_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_16_ff <= lut_16_out;
    end
end

assign out_data[16] = lut_16_ff;




// LUT : 17

wire lut_17_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011100110001111111111111011100010001000000001111011101010001),
            .DEVICE(DEVICE)
        )
    i_lut_17
        (
            .in_data({
                         in_data[304],
                         in_data[221],
                         in_data[182],
                         in_data[34],
                         in_data[319],
                         in_data[77]
                    }),
            .out_data(lut_17_out)
        );

reg   lut_17_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_17_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_17_ff <= lut_17_out;
    end
end

assign out_data[17] = lut_17_ff;




// LUT : 18

wire lut_18_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100111111011011110010111111101111111111111111111111111111111111),
            .DEVICE(DEVICE)
        )
    i_lut_18
        (
            .in_data({
                         in_data[152],
                         in_data[216],
                         in_data[33],
                         in_data[167],
                         in_data[291],
                         in_data[339]
                    }),
            .out_data(lut_18_out)
        );

reg   lut_18_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_18_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_18_ff <= lut_18_out;
    end
end

assign out_data[18] = lut_18_ff;




// LUT : 19

wire lut_19_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000010001110101011101110111100000000000010000000101010001110),
            .DEVICE(DEVICE)
        )
    i_lut_19
        (
            .in_data({
                         in_data[74],
                         in_data[45],
                         in_data[315],
                         in_data[4],
                         in_data[220],
                         in_data[166]
                    }),
            .out_data(lut_19_out)
        );

reg   lut_19_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_19_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_19_ff <= lut_19_out;
    end
end

assign out_data[19] = lut_19_ff;




// LUT : 20

wire lut_20_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100001000000000010000000000000011001110010010101100101001000000),
            .DEVICE(DEVICE)
        )
    i_lut_20
        (
            .in_data({
                         in_data[64],
                         in_data[266],
                         in_data[262],
                         in_data[312],
                         in_data[172],
                         in_data[21]
                    }),
            .out_data(lut_20_out)
        );

reg   lut_20_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_20_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_20_ff <= lut_20_out;
    end
end

assign out_data[20] = lut_20_ff;




// LUT : 21

wire lut_21_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110111110100010101000000010000011111111001000101011001110100000),
            .DEVICE(DEVICE)
        )
    i_lut_21
        (
            .in_data({
                         in_data[54],
                         in_data[311],
                         in_data[211],
                         in_data[51],
                         in_data[26],
                         in_data[208]
                    }),
            .out_data(lut_21_out)
        );

reg   lut_21_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_21_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_21_ff <= lut_21_out;
    end
end

assign out_data[21] = lut_21_ff;




// LUT : 22

wire lut_22_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000011000101110011001100110000000000010101010000000001000101),
            .DEVICE(DEVICE)
        )
    i_lut_22
        (
            .in_data({
                         in_data[43],
                         in_data[107],
                         in_data[1],
                         in_data[52],
                         in_data[332],
                         in_data[118]
                    }),
            .out_data(lut_22_out)
        );

reg   lut_22_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_22_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_22_ff <= lut_22_out;
    end
end

assign out_data[22] = lut_22_ff;




// LUT : 23

wire lut_23_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000101110100011100010000000000110001011101110111000100010000),
            .DEVICE(DEVICE)
        )
    i_lut_23
        (
            .in_data({
                         in_data[202],
                         in_data[188],
                         in_data[195],
                         in_data[335],
                         in_data[49],
                         in_data[35]
                    }),
            .out_data(lut_23_out)
        );

reg   lut_23_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_23_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_23_ff <= lut_23_out;
    end
end

assign out_data[23] = lut_23_ff;




// LUT : 24

wire lut_24_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100000110000111111111111111011111011001100001111101110110010),
            .DEVICE(DEVICE)
        )
    i_lut_24
        (
            .in_data({
                         in_data[17],
                         in_data[155],
                         in_data[270],
                         in_data[241],
                         in_data[149],
                         in_data[269]
                    }),
            .out_data(lut_24_out)
        );

reg   lut_24_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_24_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_24_ff <= lut_24_out;
    end
end

assign out_data[24] = lut_24_ff;




// LUT : 25

wire lut_25_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001100110011001100110001000100110011010101010001001100000101),
            .DEVICE(DEVICE)
        )
    i_lut_25
        (
            .in_data({
                         in_data[63],
                         in_data[69],
                         in_data[248],
                         in_data[142],
                         in_data[176],
                         in_data[357]
                    }),
            .out_data(lut_25_out)
        );

reg   lut_25_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_25_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_25_ff <= lut_25_out;
    end
end

assign out_data[25] = lut_25_ff;




// LUT : 26

wire lut_26_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111111111111101110101011111110111010111111111),
            .DEVICE(DEVICE)
        )
    i_lut_26
        (
            .in_data({
                         in_data[231],
                         in_data[236],
                         in_data[324],
                         in_data[11],
                         in_data[179],
                         in_data[131]
                    }),
            .out_data(lut_26_out)
        );

reg   lut_26_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_26_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_26_ff <= lut_26_out;
    end
end

assign out_data[26] = lut_26_ff;




// LUT : 27

wire lut_27_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011001000000000101100110011000010110010001100001111101111110010),
            .DEVICE(DEVICE)
        )
    i_lut_27
        (
            .in_data({
                         in_data[16],
                         in_data[164],
                         in_data[256],
                         in_data[223],
                         in_data[122],
                         in_data[86]
                    }),
            .out_data(lut_27_out)
        );

reg   lut_27_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_27_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_27_ff <= lut_27_out;
    end
end

assign out_data[27] = lut_27_ff;




// LUT : 28

wire lut_28_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110011011111000001000100110111011101111111110000010101001111),
            .DEVICE(DEVICE)
        )
    i_lut_28
        (
            .in_data({
                         in_data[80],
                         in_data[346],
                         in_data[84],
                         in_data[244],
                         in_data[2],
                         in_data[283]
                    }),
            .out_data(lut_28_out)
        );

reg   lut_28_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_28_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_28_ff <= lut_28_out;
    end
end

assign out_data[28] = lut_28_ff;




// LUT : 29

wire lut_29_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010001000100010101000100010000010101011001100111111101110110010),
            .DEVICE(DEVICE)
        )
    i_lut_29
        (
            .in_data({
                         in_data[264],
                         in_data[130],
                         in_data[186],
                         in_data[249],
                         in_data[42],
                         in_data[331]
                    }),
            .out_data(lut_29_out)
        );

reg   lut_29_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_29_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_29_ff <= lut_29_out;
    end
end

assign out_data[29] = lut_29_ff;




// LUT : 30

wire lut_30_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000000000000000000001010001111101010000000001000000),
            .DEVICE(DEVICE)
        )
    i_lut_30
        (
            .in_data({
                         in_data[286],
                         in_data[99],
                         in_data[284],
                         in_data[333],
                         in_data[151],
                         in_data[321]
                    }),
            .out_data(lut_30_out)
        );

reg   lut_30_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_30_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_30_ff <= lut_30_out;
    end
end

assign out_data[30] = lut_30_ff;




// LUT : 31

wire lut_31_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0011000011111111000000000111000111110111111111110111000111110111),
            .DEVICE(DEVICE)
        )
    i_lut_31
        (
            .in_data({
                         in_data[228],
                         in_data[67],
                         in_data[160],
                         in_data[3],
                         in_data[189],
                         in_data[243]
                    }),
            .out_data(lut_31_out)
        );

reg   lut_31_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_31_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_31_ff <= lut_31_out;
    end
end

assign out_data[31] = lut_31_ff;




// LUT : 32

wire lut_32_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001010100000001000000010000010110011101000001011001000100000),
            .DEVICE(DEVICE)
        )
    i_lut_32
        (
            .in_data({
                         in_data[60],
                         in_data[62],
                         in_data[294],
                         in_data[198],
                         in_data[229],
                         in_data[309]
                    }),
            .out_data(lut_32_out)
        );

reg   lut_32_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_32_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_32_ff <= lut_32_out;
    end
end

assign out_data[32] = lut_32_ff;




// LUT : 33

wire lut_33_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111101111111011101110001010101111111000011110111011100000111),
            .DEVICE(DEVICE)
        )
    i_lut_33
        (
            .in_data({
                         in_data[214],
                         in_data[100],
                         in_data[318],
                         in_data[207],
                         in_data[204],
                         in_data[39]
                    }),
            .out_data(lut_33_out)
        );

reg   lut_33_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_33_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_33_ff <= lut_33_out;
    end
end

assign out_data[33] = lut_33_ff;




// LUT : 34

wire lut_34_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111000101111101010100000111011101111111111111010111000101111),
            .DEVICE(DEVICE)
        )
    i_lut_34
        (
            .in_data({
                         in_data[292],
                         in_data[279],
                         in_data[76],
                         in_data[81],
                         in_data[197],
                         in_data[113]
                    }),
            .out_data(lut_34_out)
        );

reg   lut_34_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_34_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_34_ff <= lut_34_out;
    end
end

assign out_data[34] = lut_34_ff;




// LUT : 35

wire lut_35_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000011010101110100001111110100000000000000000000000011010100),
            .DEVICE(DEVICE)
        )
    i_lut_35
        (
            .in_data({
                         in_data[190],
                         in_data[14],
                         in_data[209],
                         in_data[177],
                         in_data[92],
                         in_data[314]
                    }),
            .out_data(lut_35_out)
        );

reg   lut_35_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_35_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_35_ff <= lut_35_out;
    end
end

assign out_data[35] = lut_35_ff;




// LUT : 36

wire lut_36_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0101010101010111000000000011000101010111011101110101001101110111),
            .DEVICE(DEVICE)
        )
    i_lut_36
        (
            .in_data({
                         in_data[240],
                         in_data[27],
                         in_data[290],
                         in_data[136],
                         in_data[287],
                         in_data[273]
                    }),
            .out_data(lut_36_out)
        );

reg   lut_36_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_36_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_36_ff <= lut_36_out;
    end
end

assign out_data[36] = lut_36_ff;




// LUT : 37

wire lut_37_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000010101010001000111110001001100001111011101110001),
            .DEVICE(DEVICE)
        )
    i_lut_37
        (
            .in_data({
                         in_data[22],
                         in_data[46],
                         in_data[102],
                         in_data[323],
                         in_data[351],
                         in_data[134]
                    }),
            .out_data(lut_37_out)
        );

reg   lut_37_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_37_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_37_ff <= lut_37_out;
    end
end

assign out_data[37] = lut_37_ff;




// LUT : 38

wire lut_38_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111010111111111011100011111001101110001111111110001000001110011),
            .DEVICE(DEVICE)
        )
    i_lut_38
        (
            .in_data({
                         in_data[119],
                         in_data[251],
                         in_data[169],
                         in_data[183],
                         in_data[162],
                         in_data[108]
                    }),
            .out_data(lut_38_out)
        );

reg   lut_38_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_38_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_38_ff <= lut_38_out;
    end
end

assign out_data[38] = lut_38_ff;




// LUT : 39

wire lut_39_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000001110000000100001111001101010000111100110111000111110111),
            .DEVICE(DEVICE)
        )
    i_lut_39
        (
            .in_data({
                         in_data[253],
                         in_data[215],
                         in_data[114],
                         in_data[28],
                         in_data[336],
                         in_data[328]
                    }),
            .out_data(lut_39_out)
        );

reg   lut_39_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_39_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_39_ff <= lut_39_out;
    end
end

assign out_data[39] = lut_39_ff;




// LUT : 40

wire lut_40_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111101110110010001100110010001011111111111100111011101110110011),
            .DEVICE(DEVICE)
        )
    i_lut_40
        (
            .in_data({
                         in_data[75],
                         in_data[173],
                         in_data[326],
                         in_data[127],
                         in_data[5],
                         in_data[25]
                    }),
            .out_data(lut_40_out)
        );

reg   lut_40_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_40_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_40_ff <= lut_40_out;
    end
end

assign out_data[40] = lut_40_ff;




// LUT : 41

wire lut_41_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010100010001000101110001010100111111011100010011111101111111),
            .DEVICE(DEVICE)
        )
    i_lut_41
        (
            .in_data({
                         in_data[210],
                         in_data[68],
                         in_data[225],
                         in_data[12],
                         in_data[345],
                         in_data[174]
                    }),
            .out_data(lut_41_out)
        );

reg   lut_41_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_41_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_41_ff <= lut_41_out;
    end
end

assign out_data[41] = lut_41_ff;




// LUT : 42

wire lut_42_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100000001000100011100000100000001110000010001000111000001110),
            .DEVICE(DEVICE)
        )
    i_lut_42
        (
            .in_data({
                         in_data[238],
                         in_data[139],
                         in_data[93],
                         in_data[175],
                         in_data[89],
                         in_data[230]
                    }),
            .out_data(lut_42_out)
        );

reg   lut_42_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_42_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_42_ff <= lut_42_out;
    end
end

assign out_data[42] = lut_42_ff;




// LUT : 43

wire lut_43_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1011000000100000001000000000000010111010001100100010000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_43
        (
            .in_data({
                         in_data[271],
                         in_data[138],
                         in_data[105],
                         in_data[307],
                         in_data[66],
                         in_data[91]
                    }),
            .out_data(lut_43_out)
        );

reg   lut_43_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_43_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_43_ff <= lut_43_out;
    end
end

assign out_data[43] = lut_43_ff;




// LUT : 44

wire lut_44_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111001001010110011101110011100011111111111111111011101111011111),
            .DEVICE(DEVICE)
        )
    i_lut_44
        (
            .in_data({
                         in_data[150],
                         in_data[90],
                         in_data[301],
                         in_data[233],
                         in_data[95],
                         in_data[137]
                    }),
            .out_data(lut_44_out)
        );

reg   lut_44_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_44_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_44_ff <= lut_44_out;
    end
end

assign out_data[44] = lut_44_ff;




// LUT : 45

wire lut_45_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101000111111000000000010101000000000001010110000000000001010),
            .DEVICE(DEVICE)
        )
    i_lut_45
        (
            .in_data({
                         in_data[260],
                         in_data[59],
                         in_data[145],
                         in_data[308],
                         in_data[299],
                         in_data[13]
                    }),
            .out_data(lut_45_out)
        );

reg   lut_45_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_45_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_45_ff <= lut_45_out;
    end
end

assign out_data[45] = lut_45_ff;




// LUT : 46

wire lut_46_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0100110111001101110011011100110100000100000011000100010011001101),
            .DEVICE(DEVICE)
        )
    i_lut_46
        (
            .in_data({
                         in_data[226],
                         in_data[170],
                         in_data[250],
                         in_data[354],
                         in_data[261],
                         in_data[121]
                    }),
            .out_data(lut_46_out)
        );

reg   lut_46_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_46_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_46_ff <= lut_46_out;
    end
end

assign out_data[46] = lut_46_ff;




// LUT : 47

wire lut_47_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111100010100000101100000010000011111011001100001011101000110000),
            .DEVICE(DEVICE)
        )
    i_lut_47
        (
            .in_data({
                         in_data[297],
                         in_data[70],
                         in_data[285],
                         in_data[288],
                         in_data[180],
                         in_data[83]
                    }),
            .out_data(lut_47_out)
        );

reg   lut_47_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_47_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_47_ff <= lut_47_out;
    end
end

assign out_data[47] = lut_47_ff;




// LUT : 48

wire lut_48_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0010101000001000101010110010101000001010000010000010101000001010),
            .DEVICE(DEVICE)
        )
    i_lut_48
        (
            .in_data({
                         in_data[55],
                         in_data[184],
                         in_data[117],
                         in_data[303],
                         in_data[245],
                         in_data[349]
                    }),
            .out_data(lut_48_out)
        );

reg   lut_48_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_48_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_48_ff <= lut_48_out;
    end
end

assign out_data[48] = lut_48_ff;




// LUT : 49

wire lut_49_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000100010011000100010111111100000000000000110000000000000011),
            .DEVICE(DEVICE)
        )
    i_lut_49
        (
            .in_data({
                         in_data[246],
                         in_data[161],
                         in_data[163],
                         in_data[50],
                         in_data[140],
                         in_data[56]
                    }),
            .out_data(lut_49_out)
        );

reg   lut_49_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_49_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_49_ff <= lut_49_out;
    end
end

assign out_data[49] = lut_49_ff;




// LUT : 50

wire lut_50_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111111111111111111101111111011111110111111001111111011111100),
            .DEVICE(DEVICE)
        )
    i_lut_50
        (
            .in_data({
                         in_data[306],
                         in_data[356],
                         in_data[277],
                         in_data[268],
                         in_data[358],
                         in_data[109]
                    }),
            .out_data(lut_50_out)
        );

reg   lut_50_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_50_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_50_ff <= lut_50_out;
    end
end

assign out_data[50] = lut_50_ff;




// LUT : 51

wire lut_51_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111110000000100000000000000100001111000001010001010100000101),
            .DEVICE(DEVICE)
        )
    i_lut_51
        (
            .in_data({
                         in_data[219],
                         in_data[213],
                         in_data[305],
                         in_data[9],
                         in_data[143],
                         in_data[199]
                    }),
            .out_data(lut_51_out)
        );

reg   lut_51_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_51_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_51_ff <= lut_51_out;
    end
end

assign out_data[51] = lut_51_ff;




// LUT : 52

wire lut_52_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000101100000010000000000000000000000010000000100000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_52
        (
            .in_data({
                         in_data[165],
                         in_data[154],
                         in_data[126],
                         in_data[87],
                         in_data[31],
                         in_data[342]
                    }),
            .out_data(lut_52_out)
        );

reg   lut_52_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_52_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_52_ff <= lut_52_out;
    end
end

assign out_data[52] = lut_52_ff;




// LUT : 53

wire lut_53_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000100000000000100011100000100000000000000000001000111000001000),
            .DEVICE(DEVICE)
        )
    i_lut_53
        (
            .in_data({
                         in_data[7],
                         in_data[153],
                         in_data[300],
                         in_data[212],
                         in_data[281],
                         in_data[192]
                    }),
            .out_data(lut_53_out)
        );

reg   lut_53_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_53_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_53_ff <= lut_53_out;
    end
end

assign out_data[53] = lut_53_ff;




// LUT : 54

wire lut_54_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000000000000000010000000000000001000000000000001101010111000000),
            .DEVICE(DEVICE)
        )
    i_lut_54
        (
            .in_data({
                         in_data[23],
                         in_data[313],
                         in_data[239],
                         in_data[6],
                         in_data[110],
                         in_data[29]
                    }),
            .out_data(lut_54_out)
        );

reg   lut_54_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_54_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_54_ff <= lut_54_out;
    end
end

assign out_data[54] = lut_54_ff;




// LUT : 55

wire lut_55_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111010111111111110001001101010111111101111111111101110111111111),
            .DEVICE(DEVICE)
        )
    i_lut_55
        (
            .in_data({
                         in_data[255],
                         in_data[15],
                         in_data[227],
                         in_data[85],
                         in_data[18],
                         in_data[196]
                    }),
            .out_data(lut_55_out)
        );

reg   lut_55_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_55_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_55_ff <= lut_55_out;
    end
end

assign out_data[55] = lut_55_ff;




// LUT : 56

wire lut_56_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1100110100001100010011000000010001001100000001000000010000000100),
            .DEVICE(DEVICE)
        )
    i_lut_56
        (
            .in_data({
                         in_data[38],
                         in_data[217],
                         in_data[106],
                         in_data[103],
                         in_data[57],
                         in_data[24]
                    }),
            .out_data(lut_56_out)
        );

reg   lut_56_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_56_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_56_ff <= lut_56_out;
    end
end

assign out_data[56] = lut_56_ff;




// LUT : 57

wire lut_57_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0001000011110101000100000101010000110011111101110000000001110011),
            .DEVICE(DEVICE)
        )
    i_lut_57
        (
            .in_data({
                         in_data[237],
                         in_data[146],
                         in_data[156],
                         in_data[242],
                         in_data[282],
                         in_data[257]
                    }),
            .out_data(lut_57_out)
        );

reg   lut_57_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_57_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_57_ff <= lut_57_out;
    end
end

assign out_data[57] = lut_57_ff;




// LUT : 58

wire lut_58_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111000111110111000100000111000111110111111111110011000011110111),
            .DEVICE(DEVICE)
        )
    i_lut_58
        (
            .in_data({
                         in_data[185],
                         in_data[158],
                         in_data[350],
                         in_data[343],
                         in_data[325],
                         in_data[88]
                    }),
            .out_data(lut_58_out)
        );

reg   lut_58_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_58_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_58_ff <= lut_58_out;
    end
end

assign out_data[58] = lut_58_ff;




// LUT : 59

wire lut_59_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0000010100000001011111110011001100000001000000000001010100000001),
            .DEVICE(DEVICE)
        )
    i_lut_59
        (
            .in_data({
                         in_data[72],
                         in_data[295],
                         in_data[258],
                         in_data[187],
                         in_data[348],
                         in_data[201]
                    }),
            .out_data(lut_59_out)
        );

reg   lut_59_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_59_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_59_ff <= lut_59_out;
    end
end

assign out_data[59] = lut_59_ff;



endmodule



module MnistStochasticLut6Mlp_sub3
        #(
            parameter DEVICE = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [59:0]  in_data,
            output wire [9:0]  out_data
        );


// LUT : 0

wire lut_0_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b0111111100110111000101110000000111111111111111110111111100010111),
            .DEVICE(DEVICE)
        )
    i_lut_0
        (
            .in_data({
                         in_data[33],
                         in_data[52],
                         in_data[32],
                         in_data[27],
                         in_data[17],
                         in_data[8]
                    }),
            .out_data(lut_0_out)
        );

reg   lut_0_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_0_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_0_ff <= lut_0_out;
    end
end

assign out_data[0] = lut_0_ff;




// LUT : 1

wire lut_1_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111111011101000100000001000000011111000100000001000000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_1
        (
            .in_data({
                         in_data[20],
                         in_data[53],
                         in_data[14],
                         in_data[26],
                         in_data[25],
                         in_data[51]
                    }),
            .out_data(lut_1_out)
        );

reg   lut_1_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_1_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_1_ff <= lut_1_out;
    end
end

assign out_data[1] = lut_1_ff;




// LUT : 2

wire lut_2_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1110100010000000111110001100000011111010111010001111111011111000),
            .DEVICE(DEVICE)
        )
    i_lut_2
        (
            .in_data({
                         in_data[57],
                         in_data[16],
                         in_data[47],
                         in_data[10],
                         in_data[3],
                         in_data[24]
                    }),
            .out_data(lut_2_out)
        );

reg   lut_2_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_2_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_2_ff <= lut_2_out;
    end
end

assign out_data[2] = lut_2_ff;




// LUT : 3

wire lut_3_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1010111111111111000010101010111100001010101011110000000000001010),
            .DEVICE(DEVICE)
        )
    i_lut_3
        (
            .in_data({
                         in_data[37],
                         in_data[21],
                         in_data[58],
                         in_data[22],
                         in_data[44],
                         in_data[19]
                    }),
            .out_data(lut_3_out)
        );

reg   lut_3_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_3_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_3_ff <= lut_3_out;
    end
end

assign out_data[3] = lut_3_ff;




// LUT : 4

wire lut_4_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011101110001111111111111011101110001000000001111011101110001),
            .DEVICE(DEVICE)
        )
    i_lut_4
        (
            .in_data({
                         in_data[45],
                         in_data[31],
                         in_data[48],
                         in_data[9],
                         in_data[7],
                         in_data[15]
                    }),
            .out_data(lut_4_out)
        );

reg   lut_4_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_4_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_4_ff <= lut_4_out;
    end
end

assign out_data[4] = lut_4_ff;




// LUT : 5

wire lut_5_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110101011101111111111101111101001101000001001101111101001101),
            .DEVICE(DEVICE)
        )
    i_lut_5
        (
            .in_data({
                         in_data[0],
                         in_data[28],
                         in_data[30],
                         in_data[34],
                         in_data[2],
                         in_data[41]
                    }),
            .out_data(lut_5_out)
        );

reg   lut_5_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_5_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_5_ff <= lut_5_out;
    end
end

assign out_data[5] = lut_5_ff;




// LUT : 6

wire lut_6_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101110111010100110001000100000011111111110101001101110001000000),
            .DEVICE(DEVICE)
        )
    i_lut_6
        (
            .in_data({
                         in_data[18],
                         in_data[54],
                         in_data[35],
                         in_data[40],
                         in_data[1],
                         in_data[50]
                    }),
            .out_data(lut_6_out)
        );

reg   lut_6_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_6_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_6_ff <= lut_6_out;
    end
end

assign out_data[6] = lut_6_ff;




// LUT : 7

wire lut_7_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1101010111000100111111111101110011000100000000001111110111000100),
            .DEVICE(DEVICE)
        )
    i_lut_7
        (
            .in_data({
                         in_data[46],
                         in_data[38],
                         in_data[36],
                         in_data[42],
                         in_data[6],
                         in_data[4]
                    }),
            .out_data(lut_7_out)
        );

reg   lut_7_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_7_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_7_ff <= lut_7_out;
    end
end

assign out_data[7] = lut_7_ff;




// LUT : 8

wire lut_8_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1111011101110001011100010001000001110001000100000001000000000000),
            .DEVICE(DEVICE)
        )
    i_lut_8
        (
            .in_data({
                         in_data[13],
                         in_data[29],
                         in_data[39],
                         in_data[59],
                         in_data[11],
                         in_data[23]
                    }),
            .out_data(lut_8_out)
        );

reg   lut_8_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_8_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_8_ff <= lut_8_out;
    end
end

assign out_data[8] = lut_8_ff;




// LUT : 9

wire lut_9_out;

bb_lut
        #(
            .N(6),
            .INIT(64'b1000111000001000111111111100111111101110100011101111111111101111),
            .DEVICE(DEVICE)
        )
    i_lut_9
        (
            .in_data({
                         in_data[43],
                         in_data[12],
                         in_data[49],
                         in_data[55],
                         in_data[56],
                         in_data[5]
                    }),
            .out_data(lut_9_out)
        );

reg   lut_9_ff;
always @(posedge clk) begin
    if ( reset ) begin
        lut_9_ff <= 1'b0;
    end
    else if ( cke ) begin
        lut_9_ff <= lut_9_out;
    end
end

assign out_data[9] = lut_9_ff;



endmodule

